magic
tech gf180mcuC
magscale 1 5
timestamp 1670312215
<< obsm1 >>
rect 672 855 189280 188190
<< metal2 >>
rect 3192 189600 3248 190000
rect 4816 189600 4872 190000
rect 6440 189600 6496 190000
rect 8064 189600 8120 190000
rect 9688 189600 9744 190000
rect 11312 189600 11368 190000
rect 12936 189600 12992 190000
rect 14560 189600 14616 190000
rect 16184 189600 16240 190000
rect 17808 189600 17864 190000
rect 19432 189600 19488 190000
rect 21056 189600 21112 190000
rect 22680 189600 22736 190000
rect 24304 189600 24360 190000
rect 25928 189600 25984 190000
rect 27552 189600 27608 190000
rect 29176 189600 29232 190000
rect 30800 189600 30856 190000
rect 32424 189600 32480 190000
rect 34048 189600 34104 190000
rect 35672 189600 35728 190000
rect 37296 189600 37352 190000
rect 38920 189600 38976 190000
rect 40544 189600 40600 190000
rect 42168 189600 42224 190000
rect 43792 189600 43848 190000
rect 45416 189600 45472 190000
rect 47040 189600 47096 190000
rect 48664 189600 48720 190000
rect 50288 189600 50344 190000
rect 51912 189600 51968 190000
rect 53536 189600 53592 190000
rect 55160 189600 55216 190000
rect 56784 189600 56840 190000
rect 58408 189600 58464 190000
rect 60032 189600 60088 190000
rect 61656 189600 61712 190000
rect 63280 189600 63336 190000
rect 64904 189600 64960 190000
rect 66528 189600 66584 190000
rect 68152 189600 68208 190000
rect 69776 189600 69832 190000
rect 71400 189600 71456 190000
rect 73024 189600 73080 190000
rect 74648 189600 74704 190000
rect 76272 189600 76328 190000
rect 77896 189600 77952 190000
rect 79520 189600 79576 190000
rect 81144 189600 81200 190000
rect 82768 189600 82824 190000
rect 84392 189600 84448 190000
rect 86016 189600 86072 190000
rect 87640 189600 87696 190000
rect 89264 189600 89320 190000
rect 90888 189600 90944 190000
rect 92512 189600 92568 190000
rect 94136 189600 94192 190000
rect 95760 189600 95816 190000
rect 97384 189600 97440 190000
rect 99008 189600 99064 190000
rect 100632 189600 100688 190000
rect 102256 189600 102312 190000
rect 103880 189600 103936 190000
rect 105504 189600 105560 190000
rect 107128 189600 107184 190000
rect 108752 189600 108808 190000
rect 110376 189600 110432 190000
rect 112000 189600 112056 190000
rect 113624 189600 113680 190000
rect 115248 189600 115304 190000
rect 116872 189600 116928 190000
rect 118496 189600 118552 190000
rect 120120 189600 120176 190000
rect 121744 189600 121800 190000
rect 123368 189600 123424 190000
rect 124992 189600 125048 190000
rect 126616 189600 126672 190000
rect 128240 189600 128296 190000
rect 129864 189600 129920 190000
rect 131488 189600 131544 190000
rect 133112 189600 133168 190000
rect 134736 189600 134792 190000
rect 136360 189600 136416 190000
rect 137984 189600 138040 190000
rect 139608 189600 139664 190000
rect 141232 189600 141288 190000
rect 142856 189600 142912 190000
rect 144480 189600 144536 190000
rect 146104 189600 146160 190000
rect 147728 189600 147784 190000
rect 149352 189600 149408 190000
rect 150976 189600 151032 190000
rect 152600 189600 152656 190000
rect 154224 189600 154280 190000
rect 155848 189600 155904 190000
rect 157472 189600 157528 190000
rect 159096 189600 159152 190000
rect 160720 189600 160776 190000
rect 162344 189600 162400 190000
rect 163968 189600 164024 190000
rect 165592 189600 165648 190000
rect 167216 189600 167272 190000
rect 168840 189600 168896 190000
rect 170464 189600 170520 190000
rect 172088 189600 172144 190000
rect 173712 189600 173768 190000
rect 175336 189600 175392 190000
rect 176960 189600 177016 190000
rect 178584 189600 178640 190000
rect 180208 189600 180264 190000
rect 181832 189600 181888 190000
rect 183456 189600 183512 190000
rect 185080 189600 185136 190000
rect 186704 189600 186760 190000
rect 2576 0 2632 400
rect 3192 0 3248 400
rect 3808 0 3864 400
rect 4424 0 4480 400
rect 5040 0 5096 400
rect 5656 0 5712 400
rect 6272 0 6328 400
rect 6888 0 6944 400
rect 7504 0 7560 400
rect 8120 0 8176 400
rect 8736 0 8792 400
rect 9352 0 9408 400
rect 9968 0 10024 400
rect 10584 0 10640 400
rect 11200 0 11256 400
rect 11816 0 11872 400
rect 12432 0 12488 400
rect 13048 0 13104 400
rect 13664 0 13720 400
rect 14280 0 14336 400
rect 14896 0 14952 400
rect 15512 0 15568 400
rect 16128 0 16184 400
rect 16744 0 16800 400
rect 17360 0 17416 400
rect 17976 0 18032 400
rect 18592 0 18648 400
rect 19208 0 19264 400
rect 19824 0 19880 400
rect 20440 0 20496 400
rect 21056 0 21112 400
rect 21672 0 21728 400
rect 22288 0 22344 400
rect 22904 0 22960 400
rect 23520 0 23576 400
rect 24136 0 24192 400
rect 24752 0 24808 400
rect 25368 0 25424 400
rect 25984 0 26040 400
rect 26600 0 26656 400
rect 27216 0 27272 400
rect 27832 0 27888 400
rect 28448 0 28504 400
rect 29064 0 29120 400
rect 29680 0 29736 400
rect 30296 0 30352 400
rect 30912 0 30968 400
rect 31528 0 31584 400
rect 32144 0 32200 400
rect 32760 0 32816 400
rect 33376 0 33432 400
rect 33992 0 34048 400
rect 34608 0 34664 400
rect 35224 0 35280 400
rect 35840 0 35896 400
rect 36456 0 36512 400
rect 37072 0 37128 400
rect 37688 0 37744 400
rect 38304 0 38360 400
rect 38920 0 38976 400
rect 39536 0 39592 400
rect 40152 0 40208 400
rect 40768 0 40824 400
rect 41384 0 41440 400
rect 42000 0 42056 400
rect 42616 0 42672 400
rect 43232 0 43288 400
rect 43848 0 43904 400
rect 44464 0 44520 400
rect 45080 0 45136 400
rect 45696 0 45752 400
rect 46312 0 46368 400
rect 46928 0 46984 400
rect 47544 0 47600 400
rect 48160 0 48216 400
rect 48776 0 48832 400
rect 49392 0 49448 400
rect 50008 0 50064 400
rect 50624 0 50680 400
rect 51240 0 51296 400
rect 51856 0 51912 400
rect 52472 0 52528 400
rect 53088 0 53144 400
rect 53704 0 53760 400
rect 54320 0 54376 400
rect 54936 0 54992 400
rect 55552 0 55608 400
rect 56168 0 56224 400
rect 56784 0 56840 400
rect 57400 0 57456 400
rect 58016 0 58072 400
rect 58632 0 58688 400
rect 59248 0 59304 400
rect 59864 0 59920 400
rect 60480 0 60536 400
rect 61096 0 61152 400
rect 61712 0 61768 400
rect 62328 0 62384 400
rect 62944 0 63000 400
rect 63560 0 63616 400
rect 64176 0 64232 400
rect 64792 0 64848 400
rect 65408 0 65464 400
rect 66024 0 66080 400
rect 66640 0 66696 400
rect 67256 0 67312 400
rect 67872 0 67928 400
rect 68488 0 68544 400
rect 69104 0 69160 400
rect 69720 0 69776 400
rect 70336 0 70392 400
rect 70952 0 71008 400
rect 71568 0 71624 400
rect 72184 0 72240 400
rect 72800 0 72856 400
rect 73416 0 73472 400
rect 74032 0 74088 400
rect 74648 0 74704 400
rect 75264 0 75320 400
rect 75880 0 75936 400
rect 76496 0 76552 400
rect 77112 0 77168 400
rect 77728 0 77784 400
rect 78344 0 78400 400
rect 78960 0 79016 400
rect 79576 0 79632 400
rect 80192 0 80248 400
rect 80808 0 80864 400
rect 81424 0 81480 400
rect 82040 0 82096 400
rect 82656 0 82712 400
rect 83272 0 83328 400
rect 83888 0 83944 400
rect 84504 0 84560 400
rect 85120 0 85176 400
rect 85736 0 85792 400
rect 86352 0 86408 400
rect 86968 0 87024 400
rect 87584 0 87640 400
rect 88200 0 88256 400
rect 88816 0 88872 400
rect 89432 0 89488 400
rect 90048 0 90104 400
rect 90664 0 90720 400
rect 91280 0 91336 400
rect 91896 0 91952 400
rect 92512 0 92568 400
rect 93128 0 93184 400
rect 93744 0 93800 400
rect 94360 0 94416 400
rect 94976 0 95032 400
rect 95592 0 95648 400
rect 96208 0 96264 400
rect 96824 0 96880 400
rect 97440 0 97496 400
rect 98056 0 98112 400
rect 98672 0 98728 400
rect 99288 0 99344 400
rect 99904 0 99960 400
rect 100520 0 100576 400
rect 101136 0 101192 400
rect 101752 0 101808 400
rect 102368 0 102424 400
rect 102984 0 103040 400
rect 103600 0 103656 400
rect 104216 0 104272 400
rect 104832 0 104888 400
rect 105448 0 105504 400
rect 106064 0 106120 400
rect 106680 0 106736 400
rect 107296 0 107352 400
rect 107912 0 107968 400
rect 108528 0 108584 400
rect 109144 0 109200 400
rect 109760 0 109816 400
rect 110376 0 110432 400
rect 110992 0 111048 400
rect 111608 0 111664 400
rect 112224 0 112280 400
rect 112840 0 112896 400
rect 113456 0 113512 400
rect 114072 0 114128 400
rect 114688 0 114744 400
rect 115304 0 115360 400
rect 115920 0 115976 400
rect 116536 0 116592 400
rect 117152 0 117208 400
rect 117768 0 117824 400
rect 118384 0 118440 400
rect 119000 0 119056 400
rect 119616 0 119672 400
rect 120232 0 120288 400
rect 120848 0 120904 400
rect 121464 0 121520 400
rect 122080 0 122136 400
rect 122696 0 122752 400
rect 123312 0 123368 400
rect 123928 0 123984 400
rect 124544 0 124600 400
rect 125160 0 125216 400
rect 125776 0 125832 400
rect 126392 0 126448 400
rect 127008 0 127064 400
rect 127624 0 127680 400
rect 128240 0 128296 400
rect 128856 0 128912 400
rect 129472 0 129528 400
rect 130088 0 130144 400
rect 130704 0 130760 400
rect 131320 0 131376 400
rect 131936 0 131992 400
rect 132552 0 132608 400
rect 133168 0 133224 400
rect 133784 0 133840 400
rect 134400 0 134456 400
rect 135016 0 135072 400
rect 135632 0 135688 400
rect 136248 0 136304 400
rect 136864 0 136920 400
rect 137480 0 137536 400
rect 138096 0 138152 400
rect 138712 0 138768 400
rect 139328 0 139384 400
rect 139944 0 140000 400
rect 140560 0 140616 400
rect 141176 0 141232 400
rect 141792 0 141848 400
rect 142408 0 142464 400
rect 143024 0 143080 400
rect 143640 0 143696 400
rect 144256 0 144312 400
rect 144872 0 144928 400
rect 145488 0 145544 400
rect 146104 0 146160 400
rect 146720 0 146776 400
rect 147336 0 147392 400
rect 147952 0 148008 400
rect 148568 0 148624 400
rect 149184 0 149240 400
rect 149800 0 149856 400
rect 150416 0 150472 400
rect 151032 0 151088 400
rect 151648 0 151704 400
rect 152264 0 152320 400
rect 152880 0 152936 400
rect 153496 0 153552 400
rect 154112 0 154168 400
rect 154728 0 154784 400
rect 155344 0 155400 400
rect 155960 0 156016 400
rect 156576 0 156632 400
rect 157192 0 157248 400
rect 157808 0 157864 400
rect 158424 0 158480 400
rect 159040 0 159096 400
rect 159656 0 159712 400
rect 160272 0 160328 400
rect 160888 0 160944 400
rect 161504 0 161560 400
rect 162120 0 162176 400
rect 162736 0 162792 400
rect 163352 0 163408 400
rect 163968 0 164024 400
rect 164584 0 164640 400
rect 165200 0 165256 400
rect 165816 0 165872 400
rect 166432 0 166488 400
rect 167048 0 167104 400
rect 167664 0 167720 400
rect 168280 0 168336 400
rect 168896 0 168952 400
rect 169512 0 169568 400
rect 170128 0 170184 400
rect 170744 0 170800 400
rect 171360 0 171416 400
rect 171976 0 172032 400
rect 172592 0 172648 400
rect 173208 0 173264 400
rect 173824 0 173880 400
rect 174440 0 174496 400
rect 175056 0 175112 400
rect 175672 0 175728 400
rect 176288 0 176344 400
rect 176904 0 176960 400
rect 177520 0 177576 400
rect 178136 0 178192 400
rect 178752 0 178808 400
rect 179368 0 179424 400
rect 179984 0 180040 400
rect 180600 0 180656 400
rect 181216 0 181272 400
rect 181832 0 181888 400
rect 182448 0 182504 400
rect 183064 0 183120 400
rect 183680 0 183736 400
rect 184296 0 184352 400
rect 184912 0 184968 400
rect 185528 0 185584 400
rect 186144 0 186200 400
rect 186760 0 186816 400
rect 187376 0 187432 400
<< obsm2 >>
rect 574 189570 3162 189600
rect 3278 189570 4786 189600
rect 4902 189570 6410 189600
rect 6526 189570 8034 189600
rect 8150 189570 9658 189600
rect 9774 189570 11282 189600
rect 11398 189570 12906 189600
rect 13022 189570 14530 189600
rect 14646 189570 16154 189600
rect 16270 189570 17778 189600
rect 17894 189570 19402 189600
rect 19518 189570 21026 189600
rect 21142 189570 22650 189600
rect 22766 189570 24274 189600
rect 24390 189570 25898 189600
rect 26014 189570 27522 189600
rect 27638 189570 29146 189600
rect 29262 189570 30770 189600
rect 30886 189570 32394 189600
rect 32510 189570 34018 189600
rect 34134 189570 35642 189600
rect 35758 189570 37266 189600
rect 37382 189570 38890 189600
rect 39006 189570 40514 189600
rect 40630 189570 42138 189600
rect 42254 189570 43762 189600
rect 43878 189570 45386 189600
rect 45502 189570 47010 189600
rect 47126 189570 48634 189600
rect 48750 189570 50258 189600
rect 50374 189570 51882 189600
rect 51998 189570 53506 189600
rect 53622 189570 55130 189600
rect 55246 189570 56754 189600
rect 56870 189570 58378 189600
rect 58494 189570 60002 189600
rect 60118 189570 61626 189600
rect 61742 189570 63250 189600
rect 63366 189570 64874 189600
rect 64990 189570 66498 189600
rect 66614 189570 68122 189600
rect 68238 189570 69746 189600
rect 69862 189570 71370 189600
rect 71486 189570 72994 189600
rect 73110 189570 74618 189600
rect 74734 189570 76242 189600
rect 76358 189570 77866 189600
rect 77982 189570 79490 189600
rect 79606 189570 81114 189600
rect 81230 189570 82738 189600
rect 82854 189570 84362 189600
rect 84478 189570 85986 189600
rect 86102 189570 87610 189600
rect 87726 189570 89234 189600
rect 89350 189570 90858 189600
rect 90974 189570 92482 189600
rect 92598 189570 94106 189600
rect 94222 189570 95730 189600
rect 95846 189570 97354 189600
rect 97470 189570 98978 189600
rect 99094 189570 100602 189600
rect 100718 189570 102226 189600
rect 102342 189570 103850 189600
rect 103966 189570 105474 189600
rect 105590 189570 107098 189600
rect 107214 189570 108722 189600
rect 108838 189570 110346 189600
rect 110462 189570 111970 189600
rect 112086 189570 113594 189600
rect 113710 189570 115218 189600
rect 115334 189570 116842 189600
rect 116958 189570 118466 189600
rect 118582 189570 120090 189600
rect 120206 189570 121714 189600
rect 121830 189570 123338 189600
rect 123454 189570 124962 189600
rect 125078 189570 126586 189600
rect 126702 189570 128210 189600
rect 128326 189570 129834 189600
rect 129950 189570 131458 189600
rect 131574 189570 133082 189600
rect 133198 189570 134706 189600
rect 134822 189570 136330 189600
rect 136446 189570 137954 189600
rect 138070 189570 139578 189600
rect 139694 189570 141202 189600
rect 141318 189570 142826 189600
rect 142942 189570 144450 189600
rect 144566 189570 146074 189600
rect 146190 189570 147698 189600
rect 147814 189570 149322 189600
rect 149438 189570 150946 189600
rect 151062 189570 152570 189600
rect 152686 189570 154194 189600
rect 154310 189570 155818 189600
rect 155934 189570 157442 189600
rect 157558 189570 159066 189600
rect 159182 189570 160690 189600
rect 160806 189570 162314 189600
rect 162430 189570 163938 189600
rect 164054 189570 165562 189600
rect 165678 189570 167186 189600
rect 167302 189570 168810 189600
rect 168926 189570 170434 189600
rect 170550 189570 172058 189600
rect 172174 189570 173682 189600
rect 173798 189570 175306 189600
rect 175422 189570 176930 189600
rect 177046 189570 178554 189600
rect 178670 189570 180178 189600
rect 180294 189570 181802 189600
rect 181918 189570 183426 189600
rect 183542 189570 185050 189600
rect 185166 189570 186674 189600
rect 186790 189570 187530 189600
rect 574 430 187530 189570
rect 574 350 2546 430
rect 2662 350 3162 430
rect 3278 350 3778 430
rect 3894 350 4394 430
rect 4510 350 5010 430
rect 5126 350 5626 430
rect 5742 350 6242 430
rect 6358 350 6858 430
rect 6974 350 7474 430
rect 7590 350 8090 430
rect 8206 350 8706 430
rect 8822 350 9322 430
rect 9438 350 9938 430
rect 10054 350 10554 430
rect 10670 350 11170 430
rect 11286 350 11786 430
rect 11902 350 12402 430
rect 12518 350 13018 430
rect 13134 350 13634 430
rect 13750 350 14250 430
rect 14366 350 14866 430
rect 14982 350 15482 430
rect 15598 350 16098 430
rect 16214 350 16714 430
rect 16830 350 17330 430
rect 17446 350 17946 430
rect 18062 350 18562 430
rect 18678 350 19178 430
rect 19294 350 19794 430
rect 19910 350 20410 430
rect 20526 350 21026 430
rect 21142 350 21642 430
rect 21758 350 22258 430
rect 22374 350 22874 430
rect 22990 350 23490 430
rect 23606 350 24106 430
rect 24222 350 24722 430
rect 24838 350 25338 430
rect 25454 350 25954 430
rect 26070 350 26570 430
rect 26686 350 27186 430
rect 27302 350 27802 430
rect 27918 350 28418 430
rect 28534 350 29034 430
rect 29150 350 29650 430
rect 29766 350 30266 430
rect 30382 350 30882 430
rect 30998 350 31498 430
rect 31614 350 32114 430
rect 32230 350 32730 430
rect 32846 350 33346 430
rect 33462 350 33962 430
rect 34078 350 34578 430
rect 34694 350 35194 430
rect 35310 350 35810 430
rect 35926 350 36426 430
rect 36542 350 37042 430
rect 37158 350 37658 430
rect 37774 350 38274 430
rect 38390 350 38890 430
rect 39006 350 39506 430
rect 39622 350 40122 430
rect 40238 350 40738 430
rect 40854 350 41354 430
rect 41470 350 41970 430
rect 42086 350 42586 430
rect 42702 350 43202 430
rect 43318 350 43818 430
rect 43934 350 44434 430
rect 44550 350 45050 430
rect 45166 350 45666 430
rect 45782 350 46282 430
rect 46398 350 46898 430
rect 47014 350 47514 430
rect 47630 350 48130 430
rect 48246 350 48746 430
rect 48862 350 49362 430
rect 49478 350 49978 430
rect 50094 350 50594 430
rect 50710 350 51210 430
rect 51326 350 51826 430
rect 51942 350 52442 430
rect 52558 350 53058 430
rect 53174 350 53674 430
rect 53790 350 54290 430
rect 54406 350 54906 430
rect 55022 350 55522 430
rect 55638 350 56138 430
rect 56254 350 56754 430
rect 56870 350 57370 430
rect 57486 350 57986 430
rect 58102 350 58602 430
rect 58718 350 59218 430
rect 59334 350 59834 430
rect 59950 350 60450 430
rect 60566 350 61066 430
rect 61182 350 61682 430
rect 61798 350 62298 430
rect 62414 350 62914 430
rect 63030 350 63530 430
rect 63646 350 64146 430
rect 64262 350 64762 430
rect 64878 350 65378 430
rect 65494 350 65994 430
rect 66110 350 66610 430
rect 66726 350 67226 430
rect 67342 350 67842 430
rect 67958 350 68458 430
rect 68574 350 69074 430
rect 69190 350 69690 430
rect 69806 350 70306 430
rect 70422 350 70922 430
rect 71038 350 71538 430
rect 71654 350 72154 430
rect 72270 350 72770 430
rect 72886 350 73386 430
rect 73502 350 74002 430
rect 74118 350 74618 430
rect 74734 350 75234 430
rect 75350 350 75850 430
rect 75966 350 76466 430
rect 76582 350 77082 430
rect 77198 350 77698 430
rect 77814 350 78314 430
rect 78430 350 78930 430
rect 79046 350 79546 430
rect 79662 350 80162 430
rect 80278 350 80778 430
rect 80894 350 81394 430
rect 81510 350 82010 430
rect 82126 350 82626 430
rect 82742 350 83242 430
rect 83358 350 83858 430
rect 83974 350 84474 430
rect 84590 350 85090 430
rect 85206 350 85706 430
rect 85822 350 86322 430
rect 86438 350 86938 430
rect 87054 350 87554 430
rect 87670 350 88170 430
rect 88286 350 88786 430
rect 88902 350 89402 430
rect 89518 350 90018 430
rect 90134 350 90634 430
rect 90750 350 91250 430
rect 91366 350 91866 430
rect 91982 350 92482 430
rect 92598 350 93098 430
rect 93214 350 93714 430
rect 93830 350 94330 430
rect 94446 350 94946 430
rect 95062 350 95562 430
rect 95678 350 96178 430
rect 96294 350 96794 430
rect 96910 350 97410 430
rect 97526 350 98026 430
rect 98142 350 98642 430
rect 98758 350 99258 430
rect 99374 350 99874 430
rect 99990 350 100490 430
rect 100606 350 101106 430
rect 101222 350 101722 430
rect 101838 350 102338 430
rect 102454 350 102954 430
rect 103070 350 103570 430
rect 103686 350 104186 430
rect 104302 350 104802 430
rect 104918 350 105418 430
rect 105534 350 106034 430
rect 106150 350 106650 430
rect 106766 350 107266 430
rect 107382 350 107882 430
rect 107998 350 108498 430
rect 108614 350 109114 430
rect 109230 350 109730 430
rect 109846 350 110346 430
rect 110462 350 110962 430
rect 111078 350 111578 430
rect 111694 350 112194 430
rect 112310 350 112810 430
rect 112926 350 113426 430
rect 113542 350 114042 430
rect 114158 350 114658 430
rect 114774 350 115274 430
rect 115390 350 115890 430
rect 116006 350 116506 430
rect 116622 350 117122 430
rect 117238 350 117738 430
rect 117854 350 118354 430
rect 118470 350 118970 430
rect 119086 350 119586 430
rect 119702 350 120202 430
rect 120318 350 120818 430
rect 120934 350 121434 430
rect 121550 350 122050 430
rect 122166 350 122666 430
rect 122782 350 123282 430
rect 123398 350 123898 430
rect 124014 350 124514 430
rect 124630 350 125130 430
rect 125246 350 125746 430
rect 125862 350 126362 430
rect 126478 350 126978 430
rect 127094 350 127594 430
rect 127710 350 128210 430
rect 128326 350 128826 430
rect 128942 350 129442 430
rect 129558 350 130058 430
rect 130174 350 130674 430
rect 130790 350 131290 430
rect 131406 350 131906 430
rect 132022 350 132522 430
rect 132638 350 133138 430
rect 133254 350 133754 430
rect 133870 350 134370 430
rect 134486 350 134986 430
rect 135102 350 135602 430
rect 135718 350 136218 430
rect 136334 350 136834 430
rect 136950 350 137450 430
rect 137566 350 138066 430
rect 138182 350 138682 430
rect 138798 350 139298 430
rect 139414 350 139914 430
rect 140030 350 140530 430
rect 140646 350 141146 430
rect 141262 350 141762 430
rect 141878 350 142378 430
rect 142494 350 142994 430
rect 143110 350 143610 430
rect 143726 350 144226 430
rect 144342 350 144842 430
rect 144958 350 145458 430
rect 145574 350 146074 430
rect 146190 350 146690 430
rect 146806 350 147306 430
rect 147422 350 147922 430
rect 148038 350 148538 430
rect 148654 350 149154 430
rect 149270 350 149770 430
rect 149886 350 150386 430
rect 150502 350 151002 430
rect 151118 350 151618 430
rect 151734 350 152234 430
rect 152350 350 152850 430
rect 152966 350 153466 430
rect 153582 350 154082 430
rect 154198 350 154698 430
rect 154814 350 155314 430
rect 155430 350 155930 430
rect 156046 350 156546 430
rect 156662 350 157162 430
rect 157278 350 157778 430
rect 157894 350 158394 430
rect 158510 350 159010 430
rect 159126 350 159626 430
rect 159742 350 160242 430
rect 160358 350 160858 430
rect 160974 350 161474 430
rect 161590 350 162090 430
rect 162206 350 162706 430
rect 162822 350 163322 430
rect 163438 350 163938 430
rect 164054 350 164554 430
rect 164670 350 165170 430
rect 165286 350 165786 430
rect 165902 350 166402 430
rect 166518 350 167018 430
rect 167134 350 167634 430
rect 167750 350 168250 430
rect 168366 350 168866 430
rect 168982 350 169482 430
rect 169598 350 170098 430
rect 170214 350 170714 430
rect 170830 350 171330 430
rect 171446 350 171946 430
rect 172062 350 172562 430
rect 172678 350 173178 430
rect 173294 350 173794 430
rect 173910 350 174410 430
rect 174526 350 175026 430
rect 175142 350 175642 430
rect 175758 350 176258 430
rect 176374 350 176874 430
rect 176990 350 177490 430
rect 177606 350 178106 430
rect 178222 350 178722 430
rect 178838 350 179338 430
rect 179454 350 179954 430
rect 180070 350 180570 430
rect 180686 350 181186 430
rect 181302 350 181802 430
rect 181918 350 182418 430
rect 182534 350 183034 430
rect 183150 350 183650 430
rect 183766 350 184266 430
rect 184382 350 184882 430
rect 184998 350 185498 430
rect 185614 350 186114 430
rect 186230 350 186730 430
rect 186846 350 187346 430
rect 187462 350 187530 430
<< obsm3 >>
rect 569 574 187143 188174
<< metal4 >>
rect 2224 1538 2384 188190
rect 9904 1538 10064 188190
rect 17584 1538 17744 188190
rect 25264 1538 25424 188190
rect 32944 1538 33104 188190
rect 40624 1538 40784 188190
rect 48304 1538 48464 188190
rect 55984 1538 56144 188190
rect 63664 1538 63824 188190
rect 71344 1538 71504 188190
rect 79024 1538 79184 188190
rect 86704 1538 86864 188190
rect 94384 1538 94544 188190
rect 102064 1538 102224 188190
rect 109744 1538 109904 188190
rect 117424 1538 117584 188190
rect 125104 1538 125264 188190
rect 132784 1538 132944 188190
rect 140464 1538 140624 188190
rect 148144 1538 148304 188190
rect 155824 1538 155984 188190
rect 163504 1538 163664 188190
rect 171184 1538 171344 188190
rect 178864 1538 179024 188190
rect 186544 1538 186704 188190
<< obsm4 >>
rect 1694 1508 2194 186975
rect 2414 1508 9874 186975
rect 10094 1508 17554 186975
rect 17774 1508 25234 186975
rect 25454 1508 32914 186975
rect 33134 1508 40594 186975
rect 40814 1508 48274 186975
rect 48494 1508 55954 186975
rect 56174 1508 63634 186975
rect 63854 1508 71314 186975
rect 71534 1508 78994 186975
rect 79214 1508 86674 186975
rect 86894 1508 94354 186975
rect 94574 1508 102034 186975
rect 102254 1508 109714 186975
rect 109934 1508 117394 186975
rect 117614 1508 125074 186975
rect 125294 1508 132754 186975
rect 132974 1508 140434 186975
rect 140654 1508 142786 186975
rect 1694 569 142786 1508
<< labels >>
rlabel metal2 s 3192 189600 3248 190000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 51912 189600 51968 190000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 56784 189600 56840 190000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 61656 189600 61712 190000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 66528 189600 66584 190000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 71400 189600 71456 190000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 76272 189600 76328 190000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 81144 189600 81200 190000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 86016 189600 86072 190000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 90888 189600 90944 190000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 95760 189600 95816 190000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8064 189600 8120 190000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 100632 189600 100688 190000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 105504 189600 105560 190000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 110376 189600 110432 190000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 115248 189600 115304 190000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 120120 189600 120176 190000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 124992 189600 125048 190000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 129864 189600 129920 190000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 134736 189600 134792 190000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 139608 189600 139664 190000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 144480 189600 144536 190000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 12936 189600 12992 190000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 149352 189600 149408 190000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 154224 189600 154280 190000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 159096 189600 159152 190000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 163968 189600 164024 190000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 168840 189600 168896 190000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 173712 189600 173768 190000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 178584 189600 178640 190000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 183456 189600 183512 190000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 17808 189600 17864 190000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 22680 189600 22736 190000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 27552 189600 27608 190000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 32424 189600 32480 190000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37296 189600 37352 190000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 42168 189600 42224 190000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 47040 189600 47096 190000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4816 189600 4872 190000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 53536 189600 53592 190000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 58408 189600 58464 190000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 63280 189600 63336 190000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 68152 189600 68208 190000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 73024 189600 73080 190000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 77896 189600 77952 190000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 82768 189600 82824 190000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 87640 189600 87696 190000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 92512 189600 92568 190000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 97384 189600 97440 190000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9688 189600 9744 190000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 102256 189600 102312 190000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 107128 189600 107184 190000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 112000 189600 112056 190000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 116872 189600 116928 190000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 121744 189600 121800 190000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 126616 189600 126672 190000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 131488 189600 131544 190000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 136360 189600 136416 190000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 141232 189600 141288 190000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 146104 189600 146160 190000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 14560 189600 14616 190000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 150976 189600 151032 190000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 155848 189600 155904 190000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 160720 189600 160776 190000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 165592 189600 165648 190000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 170464 189600 170520 190000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 175336 189600 175392 190000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 180208 189600 180264 190000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 185080 189600 185136 190000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 19432 189600 19488 190000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 24304 189600 24360 190000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 29176 189600 29232 190000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 34048 189600 34104 190000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 38920 189600 38976 190000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 43792 189600 43848 190000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 48664 189600 48720 190000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 6440 189600 6496 190000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 55160 189600 55216 190000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 60032 189600 60088 190000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 64904 189600 64960 190000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 69776 189600 69832 190000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 74648 189600 74704 190000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 79520 189600 79576 190000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 84392 189600 84448 190000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 89264 189600 89320 190000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 94136 189600 94192 190000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 99008 189600 99064 190000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11312 189600 11368 190000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 103880 189600 103936 190000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 108752 189600 108808 190000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 113624 189600 113680 190000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 118496 189600 118552 190000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 123368 189600 123424 190000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 128240 189600 128296 190000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 133112 189600 133168 190000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 137984 189600 138040 190000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 142856 189600 142912 190000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 147728 189600 147784 190000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 16184 189600 16240 190000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 152600 189600 152656 190000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 157472 189600 157528 190000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 162344 189600 162400 190000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 167216 189600 167272 190000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 172088 189600 172144 190000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 176960 189600 177016 190000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 181832 189600 181888 190000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 186704 189600 186760 190000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 21056 189600 21112 190000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 25928 189600 25984 190000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30800 189600 30856 190000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 35672 189600 35728 190000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 40544 189600 40600 190000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 45416 189600 45472 190000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 50288 189600 50344 190000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 186144 0 186200 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 186760 0 186816 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 187376 0 187432 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 67872 0 67928 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 86352 0 86408 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 88200 0 88256 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 90048 0 90104 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 91896 0 91952 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 95592 0 95648 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 97440 0 97496 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 99288 0 99344 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 101136 0 101192 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 102984 0 103040 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 69720 0 69776 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 104832 0 104888 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 106680 0 106736 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 110376 0 110432 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 112224 0 112280 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 114072 0 114128 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 115920 0 115976 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 117768 0 117824 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 119616 0 119672 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 121464 0 121520 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 71568 0 71624 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 123312 0 123368 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 125160 0 125216 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 127008 0 127064 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 128856 0 128912 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 130704 0 130760 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 132552 0 132608 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 134400 0 134456 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 136248 0 136304 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 139944 0 140000 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 73416 0 73472 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 141792 0 141848 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 143640 0 143696 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 145488 0 145544 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 147336 0 147392 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 149184 0 149240 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 151032 0 151088 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 152880 0 152936 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 154728 0 154784 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 156576 0 156632 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 158424 0 158480 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 75264 0 75320 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 160272 0 160328 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 162120 0 162176 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 163968 0 164024 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 165816 0 165872 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 169512 0 169568 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 171360 0 171416 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 173208 0 173264 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 175056 0 175112 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 176904 0 176960 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 77112 0 77168 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 178752 0 178808 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 180600 0 180656 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 182448 0 182504 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 184296 0 184352 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 80808 0 80864 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 82656 0 82712 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 84504 0 84560 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 68488 0 68544 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 86968 0 87024 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 88816 0 88872 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 90664 0 90720 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 92512 0 92568 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 94360 0 94416 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 96208 0 96264 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 98056 0 98112 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 99904 0 99960 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 101752 0 101808 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 103600 0 103656 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 70336 0 70392 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 105448 0 105504 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 107296 0 107352 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 109144 0 109200 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 110992 0 111048 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 112840 0 112896 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 114688 0 114744 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 116536 0 116592 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 118384 0 118440 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 120232 0 120288 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 122080 0 122136 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 72184 0 72240 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 123928 0 123984 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 125776 0 125832 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 127624 0 127680 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 129472 0 129528 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 131320 0 131376 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 133168 0 133224 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 135016 0 135072 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 136864 0 136920 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 138712 0 138768 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 140560 0 140616 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 74032 0 74088 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 142408 0 142464 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 144256 0 144312 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 146104 0 146160 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 147952 0 148008 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 149800 0 149856 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 151648 0 151704 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 153496 0 153552 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 155344 0 155400 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 157192 0 157248 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 159040 0 159096 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 75880 0 75936 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 160888 0 160944 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 162736 0 162792 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 164584 0 164640 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 166432 0 166488 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 168280 0 168336 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 170128 0 170184 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 171976 0 172032 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 173824 0 173880 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 175672 0 175728 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 177520 0 177576 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 77728 0 77784 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 179368 0 179424 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 181216 0 181272 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 183064 0 183120 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 184912 0 184968 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 79576 0 79632 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 81424 0 81480 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 83272 0 83328 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 85120 0 85176 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 69104 0 69160 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 87584 0 87640 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 89432 0 89488 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 91280 0 91336 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 93128 0 93184 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 94976 0 95032 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 96824 0 96880 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 98672 0 98728 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 100520 0 100576 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 102368 0 102424 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 104216 0 104272 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 70952 0 71008 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 106064 0 106120 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 107912 0 107968 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 109760 0 109816 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 111608 0 111664 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 113456 0 113512 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 115304 0 115360 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 117152 0 117208 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 119000 0 119056 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 120848 0 120904 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 122696 0 122752 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 124544 0 124600 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 126392 0 126448 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 128240 0 128296 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 130088 0 130144 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 131936 0 131992 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 133784 0 133840 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 135632 0 135688 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 137480 0 137536 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 139328 0 139384 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 141176 0 141232 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 74648 0 74704 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 144872 0 144928 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 146720 0 146776 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 148568 0 148624 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 150416 0 150472 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 152264 0 152320 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 154112 0 154168 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 155960 0 156016 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 157808 0 157864 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 159656 0 159712 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 76496 0 76552 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 161504 0 161560 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 163352 0 163408 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 165200 0 165256 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 167048 0 167104 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 168896 0 168952 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 170744 0 170800 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 172592 0 172648 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 174440 0 174496 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 176288 0 176344 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 178136 0 178192 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 78344 0 78400 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 179984 0 180040 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 181832 0 181888 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 183680 0 183736 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 185528 0 185584 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 80192 0 80248 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 82040 0 82096 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 85736 0 85792 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 188190 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 188190 6 vss
port 311 nsew ground bidirectional
rlabel metal2 s 2576 0 2632 400 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 3192 0 3248 400 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 6272 0 6328 400 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 27216 0 27272 400 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 29064 0 29120 400 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 30912 0 30968 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 32760 0 32816 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 36456 0 36512 400 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 40152 0 40208 400 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 42000 0 42056 400 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 43848 0 43904 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 45696 0 45752 400 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 47544 0 47600 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 51240 0 51296 400 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 53088 0 53144 400 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 54936 0 54992 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 58632 0 58688 400 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 60480 0 60536 400 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 62328 0 62384 400 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 66024 0 66080 400 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 17976 0 18032 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 21672 0 21728 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 25368 0 25424 400 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 4424 0 4480 400 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 27832 0 27888 400 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 31528 0 31584 400 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 35224 0 35280 400 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 38920 0 38976 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 42616 0 42672 400 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 9352 0 9408 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 46312 0 46368 400 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 51856 0 51912 400 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 53704 0 53760 400 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 55552 0 55608 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 57400 0 57456 400 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 61096 0 61152 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 62944 0 63000 400 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 11816 0 11872 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 64792 0 64848 400 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 66640 0 66696 400 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 14280 0 14336 400 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 16744 0 16800 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 20440 0 20496 400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 24136 0 24192 400 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 30296 0 30352 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 32144 0 32200 400 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 33992 0 34048 400 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 35840 0 35896 400 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 37688 0 37744 400 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 41384 0 41440 400 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 43232 0 43288 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 45080 0 45136 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 9968 0 10024 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 46928 0 46984 400 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 48776 0 48832 400 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 50624 0 50680 400 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 52472 0 52528 400 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 54320 0 54376 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 56168 0 56224 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 59864 0 59920 400 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 61712 0 61768 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 63560 0 63616 400 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 65408 0 65464 400 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 67256 0 67312 400 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 17360 0 17416 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 19208 0 19264 400 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 21056 0 21112 400 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 22904 0 22960 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 26600 0 26656 400 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 8120 0 8176 400 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 10584 0 10640 400 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 13048 0 13104 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 15512 0 15568 400 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 5656 0 5712 400 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 190000 190000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 71428466
string GDS_FILE /home/anish/projects/crypto-accelerator-chip-v3/openlane/user_proj/runs/22_12_06_02_13/results/signoff/user_proj.magic.gds
string GDS_START 347024
<< end >>

