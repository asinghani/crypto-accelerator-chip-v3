magic
tech gf180mcuC
magscale 1 10
timestamp 1670312990
<< metal1 >>
rect 82338 59390 82350 59442
rect 82402 59439 82414 59442
rect 83010 59439 83022 59442
rect 82402 59393 83022 59439
rect 82402 59390 82414 59393
rect 83010 59390 83022 59393
rect 83074 59390 83086 59442
rect 156258 59390 156270 59442
rect 156322 59439 156334 59442
rect 156930 59439 156942 59442
rect 156322 59393 156942 59439
rect 156322 59390 156334 59393
rect 156930 59390 156942 59393
rect 156994 59390 157006 59442
rect 211698 59390 211710 59442
rect 211762 59439 211774 59442
rect 212370 59439 212382 59442
rect 211762 59393 212382 59439
rect 211762 59390 211774 59393
rect 212370 59390 212382 59393
rect 212434 59390 212446 59442
rect 230178 59390 230190 59442
rect 230242 59439 230254 59442
rect 230850 59439 230862 59442
rect 230242 59393 230862 59439
rect 230242 59390 230254 59393
rect 230850 59390 230862 59393
rect 230914 59390 230926 59442
rect 322578 59390 322590 59442
rect 322642 59439 322654 59442
rect 323250 59439 323262 59442
rect 322642 59393 323262 59439
rect 322642 59390 322654 59393
rect 323250 59390 323262 59393
rect 323314 59390 323326 59442
rect 359538 59390 359550 59442
rect 359602 59439 359614 59442
rect 360210 59439 360222 59442
rect 359602 59393 360222 59439
rect 359602 59390 359614 59393
rect 360210 59390 360222 59393
rect 360274 59390 360286 59442
rect 378018 59390 378030 59442
rect 378082 59439 378094 59442
rect 378690 59439 378702 59442
rect 378082 59393 378702 59439
rect 378082 59390 378094 59393
rect 378690 59390 378702 59393
rect 378754 59390 378766 59442
rect 396498 59390 396510 59442
rect 396562 59439 396574 59442
rect 397170 59439 397182 59442
rect 396562 59393 397182 59439
rect 396562 59390 396574 59393
rect 397170 59390 397182 59393
rect 397234 59390 397246 59442
rect 414978 59390 414990 59442
rect 415042 59439 415054 59442
rect 415650 59439 415662 59442
rect 415042 59393 415662 59439
rect 415042 59390 415054 59393
rect 415650 59390 415662 59393
rect 415714 59390 415726 59442
rect 124338 59166 124350 59218
rect 124402 59215 124414 59218
rect 124898 59215 124910 59218
rect 124402 59169 124910 59215
rect 124402 59166 124414 59169
rect 124898 59166 124910 59169
rect 124962 59166 124974 59218
rect 161298 59166 161310 59218
rect 161362 59215 161374 59218
rect 161858 59215 161870 59218
rect 161362 59169 161870 59215
rect 161362 59166 161374 59169
rect 161858 59166 161870 59169
rect 161922 59166 161934 59218
rect 225138 59166 225150 59218
rect 225202 59215 225214 59218
rect 225922 59215 225934 59218
rect 225202 59169 225934 59215
rect 225202 59166 225214 59169
rect 225922 59166 225934 59169
rect 225986 59166 225998 59218
rect 262098 59166 262110 59218
rect 262162 59215 262174 59218
rect 262882 59215 262894 59218
rect 262162 59169 262894 59215
rect 262162 59166 262174 59169
rect 262882 59166 262894 59169
rect 262946 59166 262958 59218
rect 299058 59166 299070 59218
rect 299122 59215 299134 59218
rect 299842 59215 299854 59218
rect 299122 59169 299854 59215
rect 299122 59166 299134 59169
rect 299842 59166 299854 59169
rect 299906 59166 299918 59218
rect 317538 59166 317550 59218
rect 317602 59215 317614 59218
rect 318322 59215 318334 59218
rect 317602 59169 318334 59215
rect 317602 59166 317614 59169
rect 318322 59166 318334 59169
rect 318386 59166 318398 59218
rect 336018 59166 336030 59218
rect 336082 59215 336094 59218
rect 336802 59215 336814 59218
rect 336082 59169 336814 59215
rect 336082 59166 336094 59169
rect 336802 59166 336814 59169
rect 336866 59166 336878 59218
rect 354498 59166 354510 59218
rect 354562 59215 354574 59218
rect 355282 59215 355294 59218
rect 354562 59169 355294 59215
rect 354562 59166 354574 59169
rect 355282 59166 355294 59169
rect 355346 59166 355358 59218
rect 372978 59166 372990 59218
rect 373042 59215 373054 59218
rect 373762 59215 373774 59218
rect 373042 59169 373774 59215
rect 373042 59166 373054 59169
rect 373762 59166 373774 59169
rect 373826 59166 373838 59218
rect 383058 59166 383070 59218
rect 383122 59215 383134 59218
rect 383618 59215 383630 59218
rect 383122 59169 383630 59215
rect 383122 59166 383134 59169
rect 383618 59166 383630 59169
rect 383682 59166 383694 59218
rect 391458 59166 391470 59218
rect 391522 59215 391534 59218
rect 392242 59215 392254 59218
rect 391522 59169 392254 59215
rect 391522 59166 391534 59169
rect 392242 59166 392254 59169
rect 392306 59166 392318 59218
rect 401538 59166 401550 59218
rect 401602 59215 401614 59218
rect 402098 59215 402110 59218
rect 401602 59169 402110 59215
rect 401602 59166 401614 59169
rect 402098 59166 402110 59169
rect 402162 59166 402174 59218
rect 151218 59054 151230 59106
rect 151282 59103 151294 59106
rect 152002 59103 152014 59106
rect 151282 59057 152014 59103
rect 151282 59054 151294 59057
rect 152002 59054 152014 59057
rect 152066 59054 152078 59106
rect 409938 59054 409950 59106
rect 410002 59103 410014 59106
rect 410722 59103 410734 59106
rect 410002 59057 410734 59103
rect 410002 59054 410014 59057
rect 410722 59054 410734 59057
rect 410786 59054 410798 59106
rect 68898 58942 68910 58994
rect 68962 58991 68974 58994
rect 69458 58991 69470 58994
rect 68962 58945 69470 58991
rect 68962 58942 68974 58945
rect 69458 58942 69470 58945
rect 69522 58942 69534 58994
rect 198258 58942 198270 58994
rect 198322 58991 198334 58994
rect 198818 58991 198830 58994
rect 198322 58945 198830 58991
rect 198322 58942 198334 58945
rect 198818 58942 198830 58945
rect 198882 58942 198894 58994
<< via1 >>
rect 82350 59390 82402 59442
rect 83022 59390 83074 59442
rect 156270 59390 156322 59442
rect 156942 59390 156994 59442
rect 211710 59390 211762 59442
rect 212382 59390 212434 59442
rect 230190 59390 230242 59442
rect 230862 59390 230914 59442
rect 322590 59390 322642 59442
rect 323262 59390 323314 59442
rect 359550 59390 359602 59442
rect 360222 59390 360274 59442
rect 378030 59390 378082 59442
rect 378702 59390 378754 59442
rect 396510 59390 396562 59442
rect 397182 59390 397234 59442
rect 414990 59390 415042 59442
rect 415662 59390 415714 59442
rect 124350 59166 124402 59218
rect 124910 59166 124962 59218
rect 161310 59166 161362 59218
rect 161870 59166 161922 59218
rect 225150 59166 225202 59218
rect 225934 59166 225986 59218
rect 262110 59166 262162 59218
rect 262894 59166 262946 59218
rect 299070 59166 299122 59218
rect 299854 59166 299906 59218
rect 317550 59166 317602 59218
rect 318334 59166 318386 59218
rect 336030 59166 336082 59218
rect 336814 59166 336866 59218
rect 354510 59166 354562 59218
rect 355294 59166 355346 59218
rect 372990 59166 373042 59218
rect 373774 59166 373826 59218
rect 383070 59166 383122 59218
rect 383630 59166 383682 59218
rect 391470 59166 391522 59218
rect 392254 59166 392306 59218
rect 401550 59166 401602 59218
rect 402110 59166 402162 59218
rect 151230 59054 151282 59106
rect 152014 59054 152066 59106
rect 409950 59054 410002 59106
rect 410734 59054 410786 59106
rect 68910 58942 68962 58994
rect 69470 58942 69522 58994
rect 198270 58942 198322 58994
rect 198830 58942 198882 58994
<< metal2 >>
rect 10108 595644 10948 595700
rect 11032 595672 11256 597000
rect 5852 530740 5908 530750
rect 4172 516628 4228 516638
rect 2492 468916 2548 468926
rect 2492 107492 2548 468860
rect 4172 442820 4228 516572
rect 5852 462868 5908 530684
rect 5852 462802 5908 462812
rect 9212 463764 9268 463774
rect 4172 442754 4228 442764
rect 5852 447188 5908 447198
rect 5852 291060 5908 447132
rect 5852 290994 5908 291004
rect 9212 121716 9268 463708
rect 10108 442932 10164 595644
rect 10892 595476 10948 595644
rect 11004 595560 11256 595672
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 33096 595560 33348 595672
rect 55160 595560 55412 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 99288 595560 99540 595672
rect 11004 595476 11060 595560
rect 10892 595420 11060 595476
rect 33292 590548 33348 595560
rect 55356 593348 55412 595560
rect 55356 593282 55412 593292
rect 33292 590482 33348 590492
rect 12572 557844 12628 557854
rect 12572 459508 12628 557788
rect 14252 473844 14308 473854
rect 14252 461188 14308 473788
rect 14252 461122 14308 461132
rect 17612 472164 17668 472174
rect 12572 459442 12628 459452
rect 15932 457156 15988 457166
rect 14252 455700 14308 455710
rect 10108 442866 10164 442876
rect 12572 443716 12628 443726
rect 10892 438564 10948 438574
rect 10892 220500 10948 438508
rect 12572 332724 12628 443660
rect 14252 431844 14308 455644
rect 14252 431778 14308 431788
rect 12572 332658 12628 332668
rect 15932 304164 15988 457100
rect 15932 304098 15988 304108
rect 10892 220434 10948 220444
rect 9212 121650 9268 121660
rect 2492 107426 2548 107436
rect 17612 92484 17668 472108
rect 22652 470596 22708 470606
rect 19292 465556 19348 465566
rect 19292 317604 19348 465500
rect 19292 317538 19348 317548
rect 22652 191604 22708 470540
rect 22652 191538 22708 191548
rect 27692 467236 27748 467246
rect 27692 149604 27748 467180
rect 68908 465444 68964 465454
rect 36092 463876 36148 463886
rect 31052 452340 31108 452350
rect 29372 448868 29428 448878
rect 29372 176484 29428 448812
rect 31052 361284 31108 452284
rect 31052 361218 31108 361228
rect 32732 448756 32788 448766
rect 29372 176418 29428 176428
rect 27692 149538 27748 149548
rect 32732 134484 32788 448700
rect 32732 134418 32788 134428
rect 34412 440356 34468 440366
rect 17612 92418 17668 92428
rect 28588 56308 28644 56318
rect 4956 41188 5012 41198
rect 4956 36932 5012 41132
rect 4956 36866 5012 36876
rect 19292 36260 19348 36270
rect 15148 36148 15204 36158
rect 10108 22708 10164 22718
rect 10108 420 10164 22652
rect 13356 5908 13412 5918
rect 11228 480 11396 532
rect 13356 480 13412 5852
rect 15148 480 15204 36092
rect 17276 5012 17332 5022
rect 17276 480 17332 4956
rect 19292 5012 19348 36204
rect 27692 12740 27748 12750
rect 19292 4946 19348 4956
rect 22988 10948 23044 10958
rect 21084 4340 21140 4350
rect 19180 4228 19236 4238
rect 19180 480 19236 4172
rect 21084 480 21140 4284
rect 22988 480 23044 10892
rect 24892 5012 24948 5022
rect 24892 480 24948 4956
rect 27692 5012 27748 12684
rect 27692 4946 27748 4956
rect 26796 4900 26852 4910
rect 26796 480 26852 4844
rect 28588 480 28644 56252
rect 31948 52948 32004 52958
rect 30268 21028 30324 21038
rect 30268 11788 30324 20972
rect 30268 11732 30436 11788
rect 30380 480 30436 11732
rect 11228 476 11592 480
rect 11228 420 11284 476
rect 10108 364 11284 420
rect 11340 392 11592 476
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15148 392 15400 480
rect 15176 -960 15400 392
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 480
rect 30380 392 30632 480
rect 30408 -960 30632 392
rect 31948 420 32004 52892
rect 34412 50484 34468 440300
rect 36092 262164 36148 463820
rect 52892 453908 52948 453918
rect 44492 453684 44548 453694
rect 41132 452228 41188 452238
rect 37772 450436 37828 450446
rect 37772 275604 37828 450380
rect 37772 275538 37828 275548
rect 36092 262098 36148 262108
rect 41132 233604 41188 452172
rect 41132 233538 41188 233548
rect 44492 63924 44548 453628
rect 44604 449092 44660 449102
rect 44604 403284 44660 449036
rect 51212 448980 51268 448990
rect 44604 403218 44660 403228
rect 46172 447412 46228 447422
rect 46172 346164 46228 447356
rect 47852 445732 47908 445742
rect 47852 388164 47908 445676
rect 47852 388098 47908 388108
rect 49532 440468 49588 440478
rect 46172 346098 46228 346108
rect 49532 79044 49588 440412
rect 51212 163044 51268 448924
rect 52892 205044 52948 453852
rect 54572 450660 54628 450670
rect 54572 247044 54628 450604
rect 56252 443940 56308 443950
rect 56252 374724 56308 443884
rect 66444 443604 66500 443614
rect 60396 441924 60452 441934
rect 59612 440692 59668 440702
rect 59612 416724 59668 440636
rect 59612 416658 59668 416668
rect 56252 374658 56308 374668
rect 54572 246978 54628 246988
rect 52892 204978 52948 204988
rect 51212 162978 51268 162988
rect 49532 78978 49588 78988
rect 44492 63858 44548 63868
rect 56252 56420 56308 56430
rect 53788 54852 53844 54862
rect 36092 54740 36148 54750
rect 34412 50418 34468 50428
rect 34524 53060 34580 53070
rect 34524 4900 34580 53004
rect 34524 4834 34580 4844
rect 34412 4564 34468 4574
rect 32172 480 32340 532
rect 34412 480 34468 4508
rect 36092 4564 36148 54684
rect 36988 54628 37044 54638
rect 36092 4498 36148 4508
rect 36316 7588 36372 7598
rect 36316 480 36372 7532
rect 32172 476 32536 480
rect 32172 420 32228 476
rect 31948 364 32228 420
rect 32284 392 32536 476
rect 32312 -960 32536 392
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 36988 420 37044 54572
rect 40348 51268 40404 51278
rect 40124 5012 40180 5022
rect 37884 480 38052 532
rect 40124 480 40180 4956
rect 37884 476 38248 480
rect 37884 420 37940 476
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 36988 364 37940 420
rect 37996 392 38248 476
rect 38024 -960 38248 392
rect 39928 392 40180 480
rect 40348 420 40404 51212
rect 44492 27748 44548 27758
rect 44492 5012 44548 27692
rect 48748 26068 48804 26078
rect 47068 19348 47124 19358
rect 45388 17668 45444 17678
rect 45388 11788 45444 17612
rect 45388 11732 45668 11788
rect 44492 4946 44548 4956
rect 43932 4452 43988 4462
rect 41692 480 41860 532
rect 43932 480 43988 4396
rect 41692 476 42056 480
rect 41692 420 41748 476
rect 39928 -960 40152 392
rect 40348 364 41748 420
rect 41804 392 42056 476
rect 41832 -960 42056 392
rect 43736 392 43988 480
rect 45612 480 45668 11732
rect 45612 392 45864 480
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47068 420 47124 19292
rect 47404 480 47572 532
rect 47404 476 47768 480
rect 47404 420 47460 476
rect 47068 364 47460 420
rect 47516 392 47768 476
rect 47544 -960 47768 392
rect 48748 420 48804 26012
rect 52108 25172 52164 25182
rect 51548 4564 51604 4574
rect 49308 480 49476 532
rect 51548 480 51604 4508
rect 49308 476 49672 480
rect 49308 420 49364 476
rect 48748 364 49364 420
rect 49420 392 49672 476
rect 49448 -960 49672 392
rect 51352 392 51604 480
rect 52108 420 52164 25116
rect 53116 480 53284 532
rect 53116 476 53480 480
rect 53116 420 53172 476
rect 51352 -960 51576 392
rect 52108 364 53172 420
rect 53228 392 53480 476
rect 53256 -960 53480 392
rect 53788 420 53844 54796
rect 56252 25172 56308 56364
rect 56252 25106 56308 25116
rect 58828 44548 58884 44558
rect 58828 11788 58884 44492
rect 60396 42868 60452 441868
rect 66444 439880 66500 443548
rect 68908 439908 68964 465388
rect 76188 445284 76244 445294
rect 72940 441924 72996 441934
rect 68908 439852 69720 439908
rect 72940 439880 72996 441868
rect 76188 439880 76244 445228
rect 77308 443044 77364 595560
rect 99484 591332 99540 595560
rect 121324 595560 121576 595672
rect 142828 595644 143332 595700
rect 143416 595672 143640 597000
rect 99484 591266 99540 591276
rect 104972 591332 105028 591342
rect 97468 473844 97524 473854
rect 77308 442978 77364 442988
rect 78988 467124 79044 467134
rect 78988 439908 79044 467068
rect 94108 458724 94164 458734
rect 85708 457044 85764 457054
rect 82348 447076 82404 447086
rect 82348 439908 82404 447020
rect 85708 439908 85764 456988
rect 92428 452116 92484 452126
rect 89180 445508 89236 445518
rect 78988 439852 79464 439908
rect 82348 439852 82712 439908
rect 85708 439852 85960 439908
rect 89180 439880 89236 445452
rect 92428 439880 92484 452060
rect 94108 446908 94164 458668
rect 97468 446908 97524 473788
rect 104188 462084 104244 462094
rect 100828 453796 100884 453806
rect 100828 446908 100884 453740
rect 104188 446908 104244 462028
rect 104972 461412 105028 591276
rect 121324 588028 121380 595560
rect 120988 587972 121380 588028
rect 120988 474628 121044 587972
rect 120988 474562 121044 474572
rect 134428 470484 134484 470504
rect 104972 461346 105028 461356
rect 127708 462196 127764 462206
rect 117628 458948 117684 458958
rect 94108 446852 94948 446908
rect 97468 446852 98196 446908
rect 100828 446852 101444 446908
rect 104188 446852 104692 446908
rect 94892 439908 94948 446852
rect 98140 439908 98196 446852
rect 101388 439908 101444 446852
rect 104636 439908 104692 446852
rect 108668 442708 108724 442718
rect 94892 439852 95704 439908
rect 98140 439852 98952 439908
rect 101388 439852 102200 439908
rect 104636 439852 105448 439908
rect 108668 439880 108724 442652
rect 111916 441924 111972 441934
rect 111916 439880 111972 441868
rect 115164 440580 115220 440590
rect 115164 439880 115220 440524
rect 117628 439908 117684 458892
rect 124348 452004 124404 452014
rect 120988 450324 121044 450334
rect 120988 439908 121044 450268
rect 124348 439908 124404 451948
rect 127708 439908 127764 462140
rect 131068 447300 131124 447310
rect 131068 439908 131124 447244
rect 134428 439908 134484 470428
rect 142828 458052 142884 595644
rect 143276 595476 143332 595644
rect 143388 595560 143640 595672
rect 164668 595644 165396 595700
rect 165480 595672 165704 597000
rect 143388 595476 143444 595560
rect 143276 595420 143444 595476
rect 142828 457986 142884 457996
rect 142940 460404 142996 460414
rect 141148 455364 141204 455374
rect 137788 450548 137844 450558
rect 137788 439908 137844 450492
rect 117628 439852 118440 439908
rect 120988 439852 121688 439908
rect 124348 439852 124936 439908
rect 127708 439852 128184 439908
rect 131068 439852 131432 439908
rect 134428 439852 134680 439908
rect 137788 439852 137928 439908
rect 141148 439880 141204 455308
rect 142940 446908 142996 460348
rect 159628 455588 159684 455598
rect 149548 455476 149604 455486
rect 146188 450772 146244 450782
rect 146188 446908 146244 450716
rect 149548 446908 149604 455420
rect 159628 446908 159684 455532
rect 142940 446852 143668 446908
rect 146188 446852 146916 446908
rect 149548 446852 150164 446908
rect 159628 446852 159908 446908
rect 143612 439908 143668 446852
rect 146860 439908 146916 446852
rect 150108 439908 150164 446852
rect 157388 445620 157444 445630
rect 154140 443828 154196 443838
rect 143612 439852 144424 439908
rect 146860 439852 147672 439908
rect 150108 439852 150920 439908
rect 154140 439880 154196 443772
rect 157388 439880 157444 445564
rect 159852 439908 159908 446852
rect 164668 443156 164724 595644
rect 165340 595476 165396 595644
rect 165452 595560 165704 595672
rect 187544 595672 187768 597000
rect 187544 595560 187796 595672
rect 165452 595476 165508 595560
rect 165340 595420 165508 595476
rect 187740 590660 187796 595560
rect 208572 595644 209524 595700
rect 209608 595672 209832 597000
rect 187740 590594 187796 590604
rect 188972 590660 189028 590670
rect 185612 482244 185668 482254
rect 176428 468804 176484 468814
rect 170492 448644 170548 448654
rect 164668 443090 164724 443100
rect 167132 444052 167188 444062
rect 163884 440244 163940 440254
rect 159852 439852 160664 439908
rect 163884 439880 163940 440188
rect 167132 439880 167188 443996
rect 170492 442708 170548 448588
rect 170492 442642 170548 442652
rect 173068 446964 173124 446984
rect 170380 442036 170436 442046
rect 170380 439880 170436 441980
rect 173068 439908 173124 446908
rect 176428 439908 176484 468748
rect 179788 454468 179844 454478
rect 179788 439908 179844 454412
rect 183372 444164 183428 444174
rect 173068 439852 173656 439908
rect 176428 439852 176904 439908
rect 179788 439852 180152 439908
rect 183372 439880 183428 444108
rect 185612 444164 185668 482188
rect 188972 472948 189028 590604
rect 207452 588084 207508 588104
rect 194908 547764 194964 547774
rect 194012 509124 194068 509134
rect 188972 472882 189028 472892
rect 189868 495684 189924 495694
rect 185612 444098 185668 444108
rect 186620 444388 186676 444398
rect 186620 439880 186676 444332
rect 189868 439880 189924 495628
rect 191548 466228 191604 466238
rect 191548 446908 191604 466172
rect 191548 446852 192388 446908
rect 192332 439908 192388 446852
rect 194012 444388 194068 509068
rect 194908 446908 194964 547708
rect 198268 534324 198324 534334
rect 198268 446908 198324 534268
rect 201628 464548 201684 464558
rect 201628 446908 201684 464492
rect 194908 446852 195636 446908
rect 198268 446852 198884 446908
rect 201628 446852 202132 446908
rect 194012 444322 194068 444332
rect 195580 439908 195636 446852
rect 198828 439908 198884 446852
rect 202076 439908 202132 446852
rect 206108 444164 206164 444174
rect 192332 439852 193144 439908
rect 195580 439852 196392 439908
rect 198828 439852 199640 439908
rect 202076 439852 202888 439908
rect 206108 439880 206164 444108
rect 207452 444164 207508 588028
rect 208572 575428 208628 595644
rect 209468 595476 209524 595644
rect 209580 595560 209832 595672
rect 230188 595644 231588 595700
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 209580 595476 209636 595560
rect 209468 595420 209636 595476
rect 224252 593236 224308 593246
rect 208572 575362 208628 575372
rect 215068 593124 215124 593134
rect 208348 574644 208404 574654
rect 208348 446908 208404 574588
rect 212492 502404 212548 502414
rect 212492 476308 212548 502348
rect 212492 476242 212548 476252
rect 211708 467908 211764 467918
rect 211708 446908 211764 467852
rect 208348 446852 208628 446908
rect 211708 446852 211876 446908
rect 207452 444098 207508 444108
rect 208572 439908 208628 446852
rect 211820 439908 211876 446852
rect 215068 439908 215124 593068
rect 222348 443268 222404 443278
rect 219100 442708 219156 442718
rect 208572 439852 209384 439908
rect 211820 439852 212632 439908
rect 215068 439852 215880 439908
rect 219100 439880 219156 442652
rect 222348 439880 222404 443212
rect 224252 443268 224308 593180
rect 230188 464660 230244 595644
rect 231532 595476 231588 595644
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297388 595644 297780 595700
rect 297864 595672 298088 597000
rect 231644 595476 231700 595560
rect 231532 595420 231700 595476
rect 230188 464594 230244 464604
rect 231868 593460 231924 593470
rect 228508 461300 228564 461310
rect 224252 443202 224308 443212
rect 225148 457828 225204 457838
rect 225148 439908 225204 457772
rect 228508 439908 228564 461244
rect 231868 439908 231924 593404
rect 242732 590660 242788 590670
rect 238588 469588 238644 469598
rect 235228 457940 235284 457950
rect 235228 439908 235284 457884
rect 225148 439852 225624 439908
rect 228508 439852 228872 439908
rect 231868 439852 232120 439908
rect 235228 439852 235368 439908
rect 238588 439880 238644 469532
rect 241836 444164 241892 444174
rect 241836 439880 241892 444108
rect 242732 444164 242788 590604
rect 250348 503188 250404 503198
rect 246988 462980 247044 462990
rect 243628 459620 243684 459630
rect 243628 446908 243684 459564
rect 246092 458836 246148 458846
rect 246092 454580 246148 458780
rect 246092 454514 246148 454524
rect 246988 446908 247044 462924
rect 250348 446908 250404 503132
rect 253708 471268 253764 595560
rect 274652 590548 274708 590558
rect 263788 575428 263844 575438
rect 253708 471202 253764 471212
rect 260428 471268 260484 471278
rect 257068 463092 257124 463102
rect 253708 459732 253764 459742
rect 253708 446908 253764 459676
rect 257068 446908 257124 463036
rect 260428 446908 260484 471212
rect 243628 446852 244356 446908
rect 246988 446852 247604 446908
rect 250348 446852 250852 446908
rect 253708 446852 254100 446908
rect 257068 446852 257348 446908
rect 260428 446852 260596 446908
rect 242732 444098 242788 444108
rect 244300 439908 244356 446852
rect 247548 439908 247604 446852
rect 250796 439908 250852 446852
rect 254044 439908 254100 446852
rect 257292 439908 257348 446852
rect 260540 439908 260596 446852
rect 263788 439908 263844 575372
rect 270508 472948 270564 472958
rect 267148 464660 267204 464670
rect 267148 439908 267204 464604
rect 270508 439908 270564 472892
rect 273868 458052 273924 458062
rect 273868 439908 273924 457996
rect 274652 458052 274708 590492
rect 275772 588028 275828 595560
rect 275548 587972 275828 588028
rect 288988 593348 289044 593358
rect 275548 459732 275604 587972
rect 275548 459666 275604 459676
rect 280588 474628 280644 474638
rect 274652 457986 274708 457996
rect 277564 443156 277620 443166
rect 244300 439852 245112 439908
rect 247548 439852 248360 439908
rect 250796 439852 251608 439908
rect 254044 439852 254856 439908
rect 257292 439852 258104 439908
rect 260540 439852 261352 439908
rect 263788 439852 264600 439908
rect 267148 439852 267848 439908
rect 270508 439852 271096 439908
rect 273868 439852 274344 439908
rect 277564 439880 277620 443100
rect 280588 439908 280644 474572
rect 287308 461412 287364 461422
rect 284060 443044 284116 443054
rect 280588 439852 280840 439908
rect 284060 439880 284116 442988
rect 287308 439880 287364 461356
rect 288988 446908 289044 593292
rect 297388 463092 297444 595644
rect 297724 595476 297780 595644
rect 297836 595560 298088 595672
rect 319228 595644 319844 595700
rect 319928 595672 320152 597000
rect 297836 595476 297892 595560
rect 297724 595420 297892 595476
rect 303212 590548 303268 590558
rect 297388 463026 297444 463036
rect 299068 586404 299124 586414
rect 295708 458052 295764 458062
rect 295708 446908 295764 457996
rect 299068 446908 299124 586348
rect 303212 462980 303268 590492
rect 303212 462914 303268 462924
rect 305788 572964 305844 572974
rect 302428 459508 302484 459518
rect 302428 446908 302484 459452
rect 305788 446908 305844 572908
rect 308252 544404 308308 544414
rect 288988 446852 289828 446908
rect 295708 446852 296324 446908
rect 299068 446852 299572 446908
rect 302428 446852 302820 446908
rect 305788 446852 306068 446908
rect 289772 439908 289828 446852
rect 293804 442932 293860 442942
rect 289772 439852 290584 439908
rect 293804 439880 293860 442876
rect 296268 439908 296324 446852
rect 299516 439908 299572 446852
rect 302764 439908 302820 446852
rect 306012 439908 306068 446852
rect 308252 443156 308308 544348
rect 319228 503188 319284 595644
rect 319788 595476 319844 595644
rect 319900 595560 320152 595672
rect 341068 595644 341908 595700
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 319900 595476 319956 595560
rect 319788 595420 319956 595476
rect 319228 503122 319284 503132
rect 325052 487284 325108 487294
rect 319228 476308 319284 476318
rect 315868 462868 315924 462878
rect 308252 443090 308308 443100
rect 310044 443156 310100 443166
rect 296268 439852 297080 439908
rect 299516 439852 300328 439908
rect 302764 439852 303576 439908
rect 306012 439852 306824 439908
rect 310044 439880 310100 443100
rect 313292 442820 313348 442830
rect 313292 439880 313348 442764
rect 315868 439908 315924 462812
rect 319228 439908 319284 476252
rect 322588 461188 322644 461198
rect 322588 439908 322644 461132
rect 325052 448532 325108 487228
rect 341068 459620 341124 595644
rect 341852 595476 341908 595644
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 430220 595560 430472 595672
rect 451612 595644 452228 595700
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 341964 595476 342020 595560
rect 341852 595420 342020 595476
rect 364028 590548 364084 595560
rect 386092 590660 386148 595560
rect 386092 590594 386148 590604
rect 364028 590482 364084 590492
rect 393148 470596 393204 470606
rect 341068 459554 341124 459564
rect 364588 465556 364644 465566
rect 361228 457156 361284 457166
rect 332668 455700 332724 455710
rect 329308 454580 329364 454590
rect 325052 448466 325108 448476
rect 325948 448532 326004 448542
rect 325948 439908 326004 448476
rect 329308 439908 329364 454524
rect 332668 439908 332724 455644
rect 354508 452340 354564 452350
rect 344428 449092 344484 449102
rect 344428 446908 344484 449036
rect 351148 447412 351204 447422
rect 351148 446908 351204 447356
rect 354508 446908 354564 452284
rect 344428 446852 345044 446908
rect 351148 446852 351540 446908
rect 354508 446852 354788 446908
rect 342524 445732 342580 445742
rect 336028 445396 336084 445406
rect 315868 439852 316568 439908
rect 319228 439852 319816 439908
rect 322588 439852 323064 439908
rect 325948 439852 326312 439908
rect 329308 439852 329560 439908
rect 332668 439852 332808 439908
rect 336028 439880 336084 445340
rect 339276 440692 339332 440702
rect 339276 439880 339332 440636
rect 342524 439880 342580 445676
rect 344988 439908 345044 446852
rect 349020 443940 349076 443950
rect 344988 439852 345800 439908
rect 349020 439880 349076 443884
rect 351484 439908 351540 446852
rect 354732 439908 354788 446852
rect 358764 443716 358820 443726
rect 351484 439852 352296 439908
rect 354732 439852 355544 439908
rect 358764 439880 358820 443660
rect 361228 439908 361284 457100
rect 364588 439908 364644 465500
rect 371308 463876 371364 463886
rect 367948 447188 368004 447198
rect 367948 439908 368004 447132
rect 371308 439908 371364 463820
rect 386428 453908 386484 453918
rect 384748 452228 384804 452238
rect 378028 450660 378084 450670
rect 374668 450436 374724 450446
rect 374668 439908 374724 450380
rect 378028 439908 378084 450604
rect 361228 439852 362040 439908
rect 364588 439852 365288 439908
rect 367948 439852 368536 439908
rect 371308 439852 371784 439908
rect 374668 439852 375032 439908
rect 378028 439852 378280 439908
rect 384748 439880 384804 452172
rect 386428 446908 386484 453852
rect 389788 448868 389844 448878
rect 389788 446908 389844 448812
rect 393148 446908 393204 470540
rect 403228 467236 403284 467246
rect 396508 448980 396564 448990
rect 396508 446908 396564 448924
rect 399868 448756 399924 448766
rect 399868 446908 399924 448700
rect 403228 446908 403284 467180
rect 406588 463764 406644 463774
rect 406588 446908 406644 463708
rect 408268 457940 408324 595560
rect 427532 590884 427588 590894
rect 408268 457874 408324 457884
rect 409948 472164 410004 472174
rect 386428 446852 387268 446908
rect 389788 446852 390516 446908
rect 393148 446852 393764 446908
rect 396508 446852 397012 446908
rect 399868 446852 400260 446908
rect 403228 446852 403508 446908
rect 406588 446852 406756 446908
rect 387212 439908 387268 446852
rect 390460 439908 390516 446852
rect 393708 439908 393764 446852
rect 396956 439908 397012 446852
rect 400204 439908 400260 446852
rect 403452 439908 403508 446852
rect 406700 439908 406756 446852
rect 409948 439908 410004 472108
rect 427532 469588 427588 590828
rect 430220 590884 430276 595560
rect 451612 593460 451668 595644
rect 452172 595476 452228 595644
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 495628 595644 496356 595700
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 452284 595476 452340 595560
rect 452172 595420 452340 595476
rect 451612 593394 451668 593404
rect 430220 590818 430276 590828
rect 427532 469522 427588 469532
rect 454412 590548 454468 590558
rect 413308 468916 413364 468926
rect 413308 439908 413364 468860
rect 447692 462196 447748 462206
rect 444332 458948 444388 458958
rect 423388 453684 423444 453694
rect 417228 440468 417284 440478
rect 387212 439852 388024 439908
rect 390460 439852 391272 439908
rect 393708 439852 394520 439908
rect 396956 439852 397768 439908
rect 400204 439852 401016 439908
rect 403452 439852 404264 439908
rect 406700 439852 407512 439908
rect 409948 439852 410760 439908
rect 413308 439852 414008 439908
rect 417228 439880 417284 440412
rect 420476 440356 420532 440366
rect 420476 439880 420532 440300
rect 423388 439908 423444 453628
rect 442652 444052 442708 444062
rect 426972 442148 427028 442158
rect 423388 439852 423752 439908
rect 426972 439880 427028 442092
rect 440188 442148 440244 442158
rect 381500 439348 381556 439358
rect 381500 439282 381556 439292
rect 430220 439348 430276 439358
rect 430220 439282 430276 439292
rect 433468 439348 433524 439358
rect 433468 439282 433524 439292
rect 436828 438564 436884 438574
rect 63868 60060 65240 60116
rect 65548 60060 66472 60116
rect 67228 60060 67704 60116
rect 68936 60060 69076 60116
rect 60396 42802 60452 42812
rect 62972 56644 63028 56654
rect 58828 11732 58996 11788
rect 57260 4676 57316 4686
rect 55020 480 55188 532
rect 57260 480 57316 4620
rect 55020 476 55384 480
rect 55020 420 55076 476
rect 53788 364 55076 420
rect 55132 392 55384 476
rect 55160 -960 55384 392
rect 57064 392 57316 480
rect 58940 480 58996 11732
rect 62972 10948 63028 56588
rect 63868 22708 63924 60060
rect 63868 22642 63924 22652
rect 62972 10882 63028 10892
rect 63868 15988 63924 15998
rect 61068 6020 61124 6030
rect 61068 480 61124 5964
rect 62972 4788 63028 4798
rect 62972 480 63028 4732
rect 58940 392 59192 480
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 60872 392 61124 480
rect 62776 392 63028 480
rect 63868 420 63924 15932
rect 65548 5908 65604 60060
rect 67228 36148 67284 60060
rect 68908 58994 68964 59006
rect 68908 58942 68910 58994
rect 68962 58942 68964 58994
rect 67228 36082 67284 36092
rect 68012 56532 68068 56542
rect 68012 6020 68068 56476
rect 68012 5954 68068 5964
rect 65548 5842 65604 5852
rect 66780 5908 66836 5918
rect 64540 480 64708 532
rect 66780 480 66836 5852
rect 68684 4900 68740 4910
rect 68684 480 68740 4844
rect 68908 4228 68964 58942
rect 69020 36260 69076 60060
rect 69468 60060 70168 60116
rect 70588 60060 71400 60116
rect 72268 60060 72632 60116
rect 72716 60060 73864 60116
rect 73948 60060 75096 60116
rect 75628 60060 76328 60116
rect 77308 60060 77560 60116
rect 77980 60060 78792 60116
rect 78988 60060 80024 60116
rect 80668 60060 81256 60116
rect 69468 58994 69524 60060
rect 69468 58942 69470 58994
rect 69522 58942 69524 58994
rect 69468 58930 69524 58942
rect 69020 36194 69076 36204
rect 68908 4162 68964 4172
rect 69020 14308 69076 14318
rect 64540 476 64904 480
rect 64540 420 64596 476
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 63868 364 64596 420
rect 64652 392 64904 476
rect 64680 -960 64904 392
rect 66584 392 66836 480
rect 68488 392 68740 480
rect 69020 420 69076 14252
rect 70588 4340 70644 60060
rect 72268 56644 72324 60060
rect 72268 56578 72324 56588
rect 72716 12740 72772 60060
rect 73948 53060 74004 60060
rect 75628 56308 75684 60060
rect 75628 56242 75684 56252
rect 73948 52994 74004 53004
rect 76412 55524 76468 55534
rect 76412 21028 76468 55468
rect 77308 55524 77364 60060
rect 77980 58828 78036 60060
rect 77308 55458 77364 55468
rect 77420 58772 78036 58828
rect 76412 20962 76468 20972
rect 77308 53172 77364 53182
rect 72716 12674 72772 12684
rect 75628 16100 75684 16110
rect 70588 4274 70644 4284
rect 72492 12628 72548 12638
rect 70252 480 70420 532
rect 72492 480 72548 12572
rect 74396 4228 74452 4238
rect 74396 480 74452 4172
rect 70252 476 70616 480
rect 70252 420 70308 476
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 69020 364 70308 420
rect 70364 392 70616 476
rect 70392 -960 70616 392
rect 72296 392 72548 480
rect 74200 392 74452 480
rect 75628 420 75684 16044
rect 75964 480 76132 532
rect 75964 476 76328 480
rect 75964 420 76020 476
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 75628 364 76020 420
rect 76076 392 76328 476
rect 76104 -960 76328 392
rect 77308 420 77364 53116
rect 77420 52948 77476 58772
rect 78988 54740 79044 60060
rect 78988 54674 79044 54684
rect 77420 52882 77476 52892
rect 80668 7588 80724 60060
rect 82348 59442 82404 59454
rect 82348 59390 82350 59442
rect 82402 59390 82404 59442
rect 82348 27748 82404 59390
rect 82460 54628 82516 60088
rect 83020 60060 83720 60116
rect 84028 60060 84952 60116
rect 85708 60060 86184 60116
rect 83020 59442 83076 60060
rect 83020 59390 83022 59442
rect 83074 59390 83076 59442
rect 83020 59378 83076 59390
rect 82460 54562 82516 54572
rect 83132 56644 83188 56654
rect 82348 27682 82404 27692
rect 82348 21028 82404 21038
rect 80668 7522 80724 7532
rect 82012 7812 82068 7822
rect 80108 4340 80164 4350
rect 77868 480 78036 532
rect 80108 480 80164 4284
rect 82012 480 82068 7756
rect 77868 476 78232 480
rect 77868 420 77924 476
rect 77308 364 77924 420
rect 77980 392 78232 476
rect 78008 -960 78232 392
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 82348 420 82404 20972
rect 83132 5908 83188 56588
rect 84028 51268 84084 60060
rect 84028 51202 84084 51212
rect 84812 55524 84868 55534
rect 84812 17668 84868 55468
rect 84812 17602 84868 17612
rect 83132 5842 83188 5852
rect 82908 5012 82964 5022
rect 82908 4564 82964 4956
rect 82908 4498 82964 4508
rect 85708 4564 85764 60060
rect 87388 55524 87444 60088
rect 87388 55458 87444 55468
rect 87500 60060 88648 60116
rect 89068 60060 89880 60116
rect 90972 60060 91112 60116
rect 91644 60060 92344 60116
rect 92428 60060 93576 60116
rect 94108 60060 94808 60116
rect 95788 60060 96040 60116
rect 96460 60060 97272 60116
rect 97468 60060 98504 60116
rect 99148 60060 99736 60116
rect 100828 60060 100968 60116
rect 101164 60060 102200 60116
rect 102508 60060 103432 60116
rect 104188 60060 104664 60116
rect 87500 19348 87556 60060
rect 89068 26068 89124 60060
rect 90748 59444 90804 59454
rect 90748 56420 90804 59388
rect 90748 56354 90804 56364
rect 89180 55524 89236 55534
rect 89180 54852 89236 55468
rect 89180 54786 89236 54796
rect 89068 26002 89124 26012
rect 87500 19282 87556 19292
rect 89628 10948 89684 10958
rect 85708 4498 85764 4508
rect 87724 5908 87780 5918
rect 85820 4452 85876 4462
rect 83580 480 83748 532
rect 85820 480 85876 4396
rect 87724 480 87780 5852
rect 89628 480 89684 10892
rect 90972 5012 91028 60060
rect 91644 59444 91700 60060
rect 91644 59378 91700 59388
rect 91532 56756 91588 56766
rect 91532 44548 91588 56700
rect 92428 55524 92484 60060
rect 92428 55458 92484 55468
rect 91532 44482 91588 44492
rect 90972 4946 91028 4956
rect 91532 6132 91588 6142
rect 91532 480 91588 6076
rect 93436 6020 93492 6030
rect 93436 480 93492 5964
rect 94108 4676 94164 60060
rect 95788 56756 95844 60060
rect 96460 58828 96516 60060
rect 95788 56690 95844 56700
rect 95900 58772 96516 58828
rect 95900 56532 95956 58772
rect 95900 56466 95956 56476
rect 94892 56308 94948 56318
rect 94892 6132 94948 56252
rect 94892 6066 94948 6076
rect 95340 7588 95396 7598
rect 94108 4610 94164 4620
rect 95340 480 95396 7532
rect 97468 4788 97524 60060
rect 98700 56756 98756 56766
rect 98700 53172 98756 56700
rect 98700 53106 98756 53116
rect 99148 15988 99204 60060
rect 100828 56644 100884 60060
rect 101164 58828 101220 60060
rect 100828 56578 100884 56588
rect 100940 58772 101220 58828
rect 99148 15922 99204 15932
rect 99932 56532 99988 56542
rect 99932 7812 99988 56476
rect 99932 7746 99988 7756
rect 97468 4722 97524 4732
rect 99036 7700 99092 7710
rect 97244 4564 97300 4574
rect 97244 480 97300 4508
rect 99036 480 99092 7644
rect 100940 4900 100996 58772
rect 102508 14308 102564 60060
rect 102508 14242 102564 14252
rect 102732 14308 102788 14318
rect 100940 4834 100996 4844
rect 101052 4676 101108 4686
rect 101052 480 101108 4620
rect 83580 476 83944 480
rect 83580 420 83636 476
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 82348 364 83636 420
rect 83692 392 83944 476
rect 83720 -960 83944 392
rect 85624 392 85876 480
rect 87528 392 87780 480
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102732 480 102788 14252
rect 104188 12628 104244 60060
rect 104188 12562 104244 12572
rect 104412 12628 104468 12638
rect 104412 11788 104468 12572
rect 104412 11732 104692 11788
rect 104636 480 104692 11732
rect 105868 4228 105924 60088
rect 105980 60060 107128 60116
rect 107548 60060 108360 60116
rect 109452 60060 109592 60116
rect 110124 60060 110824 60116
rect 110908 60060 112056 60116
rect 112588 60060 113288 60116
rect 105980 16100 106036 60060
rect 107548 56756 107604 60060
rect 107548 56690 107604 56700
rect 109228 59444 109284 59454
rect 109228 56532 109284 59388
rect 109228 56466 109284 56476
rect 105980 16034 106036 16044
rect 107548 56420 107604 56430
rect 105868 4162 105924 4172
rect 106764 4228 106820 4238
rect 106764 480 106820 4172
rect 102732 392 102984 480
rect 104636 392 104888 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 392 106820 480
rect 107548 420 107604 56364
rect 109452 4340 109508 60060
rect 110124 59444 110180 60060
rect 110124 59378 110180 59388
rect 110012 55524 110068 55534
rect 110012 21028 110068 55468
rect 110908 55524 110964 60060
rect 110908 55458 110964 55468
rect 110012 20962 110068 20972
rect 109452 4274 109508 4284
rect 110572 6132 110628 6142
rect 108332 480 108500 532
rect 110572 480 110628 6076
rect 112588 4452 112644 60060
rect 114268 59444 114324 59454
rect 113372 55524 113428 55534
rect 113372 10948 113428 55468
rect 114268 55524 114324 59388
rect 114268 55458 114324 55468
rect 114492 55524 114548 60088
rect 115052 60060 115752 60116
rect 115948 60060 116984 60116
rect 117628 60060 118216 60116
rect 119308 60060 119448 60116
rect 119532 60060 120680 60116
rect 120988 60060 121912 60116
rect 122668 60060 123144 60116
rect 124376 60060 124516 60116
rect 115052 59444 115108 60060
rect 115052 59378 115108 59388
rect 115948 56308 116004 60060
rect 115948 56242 116004 56252
rect 114492 55458 114548 55468
rect 116060 55524 116116 55534
rect 113372 10882 113428 10892
rect 115948 15988 116004 15998
rect 115948 5908 116004 15932
rect 116060 11788 116116 55468
rect 116060 11732 116228 11788
rect 116172 5908 116228 11732
rect 117628 6020 117684 60060
rect 118412 55524 118468 55534
rect 118412 7588 118468 55468
rect 119308 55524 119364 60060
rect 119308 55458 119364 55468
rect 118412 7522 118468 7532
rect 117628 5954 117684 5964
rect 115948 5852 116116 5908
rect 112588 4386 112644 4396
rect 114380 4452 114436 4462
rect 112476 4340 112532 4350
rect 112476 480 112532 4284
rect 114380 480 114436 4396
rect 108332 476 108696 480
rect 108332 420 108388 476
rect 106568 -960 106792 392
rect 107548 364 108388 420
rect 108444 392 108696 476
rect 108472 -960 108696 392
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116060 480 116116 5852
rect 116172 5842 116228 5852
rect 118188 4788 118244 4798
rect 118188 480 118244 4732
rect 119532 4564 119588 60060
rect 119532 4498 119588 4508
rect 120092 9268 120148 9278
rect 120092 480 120148 9212
rect 120988 7700 121044 60060
rect 120988 7634 121044 7644
rect 121996 7588 122052 7598
rect 121996 480 122052 7532
rect 122668 4676 122724 60060
rect 124348 59218 124404 59230
rect 124348 59166 124350 59218
rect 124402 59166 124404 59218
rect 123452 55524 123508 55534
rect 123452 12628 123508 55468
rect 124348 55524 124404 59166
rect 124348 55458 124404 55468
rect 124460 14308 124516 60060
rect 124908 60060 125608 60116
rect 126028 60060 126840 60116
rect 127708 60060 128072 60116
rect 128492 60060 129304 60116
rect 129388 60060 130536 60116
rect 131068 60060 131768 60116
rect 132748 60060 133000 60116
rect 133420 60060 134232 60116
rect 134428 60060 135464 60116
rect 136108 60060 136696 60116
rect 137788 60060 137928 60116
rect 138124 60060 139160 60116
rect 139468 60060 140392 60116
rect 141148 60060 141624 60116
rect 142856 60060 143332 60116
rect 124908 59218 124964 60060
rect 124908 59166 124910 59218
rect 124962 59166 124964 59218
rect 124908 59154 124964 59166
rect 124460 14242 124516 14252
rect 125132 56308 125188 56318
rect 123452 12562 123508 12572
rect 122668 4610 122724 4620
rect 123900 5908 123956 5918
rect 123900 480 123956 5852
rect 125132 5908 125188 56252
rect 125132 5842 125188 5852
rect 125804 5908 125860 5918
rect 125804 480 125860 5852
rect 126028 4228 126084 60060
rect 127708 56420 127764 60060
rect 128492 58828 128548 60060
rect 127708 56354 127764 56364
rect 127820 58772 128548 58828
rect 127820 6132 127876 58772
rect 128492 56420 128548 56430
rect 128492 15988 128548 56364
rect 128492 15922 128548 15932
rect 127820 6066 127876 6076
rect 126028 4162 126084 4172
rect 127596 6020 127652 6030
rect 127596 480 127652 5964
rect 129388 4340 129444 60060
rect 131068 4452 131124 60060
rect 132748 56420 132804 60060
rect 133420 58828 133476 60060
rect 132748 56354 132804 56364
rect 132860 58772 133476 58828
rect 131852 55524 131908 55534
rect 131852 9268 131908 55468
rect 131852 9202 131908 9212
rect 131068 4386 131124 4396
rect 132636 7700 132692 7710
rect 129388 4274 129444 4284
rect 131516 3892 131572 3902
rect 129612 3444 129668 3454
rect 129612 480 129668 3388
rect 131516 480 131572 3836
rect 132636 3444 132692 7644
rect 132860 4788 132916 58772
rect 134428 55524 134484 60060
rect 134428 55458 134484 55468
rect 135212 56532 135268 56542
rect 132860 4722 132916 4732
rect 133420 5012 133476 5022
rect 132636 3378 132692 3388
rect 133420 480 133476 4956
rect 135212 5012 135268 56476
rect 135436 55524 135492 55534
rect 135436 7588 135492 55468
rect 136108 55524 136164 60060
rect 136108 55458 136164 55468
rect 136220 56420 136276 56430
rect 136220 47068 136276 56364
rect 137788 56308 137844 60060
rect 138124 58828 138180 60060
rect 137788 56242 137844 56252
rect 137900 58772 138180 58828
rect 135436 7522 135492 7532
rect 136108 47012 136276 47068
rect 135212 4946 135268 4956
rect 135324 4228 135380 4238
rect 135324 480 135380 4172
rect 116060 392 116312 480
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 392 118244 480
rect 119896 392 120148 480
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 392 129668 480
rect 131320 392 131572 480
rect 133224 392 133476 480
rect 135128 392 135380 480
rect 136108 420 136164 47012
rect 137788 7588 137844 7598
rect 137788 3892 137844 7532
rect 137900 5908 137956 58772
rect 139468 6020 139524 60060
rect 139468 5954 139524 5964
rect 140252 56644 140308 56654
rect 137900 5842 137956 5852
rect 137788 3826 137844 3836
rect 139132 5012 139188 5022
rect 136892 480 137060 532
rect 139132 480 139188 4956
rect 140252 5012 140308 56588
rect 141148 7700 141204 60060
rect 142828 59444 142884 59454
rect 142828 56532 142884 59388
rect 142828 56466 142884 56476
rect 141148 7634 141204 7644
rect 142716 8036 142772 8046
rect 140252 4946 140308 4956
rect 141036 5908 141092 5918
rect 141036 480 141092 5852
rect 142716 4228 142772 7980
rect 143276 7588 143332 60060
rect 143388 60060 144088 60116
rect 144620 60060 145320 60116
rect 146300 60060 146552 60116
rect 147084 60060 147784 60116
rect 147868 60060 149016 60116
rect 149548 60060 150248 60116
rect 151340 60060 151480 60116
rect 152012 60060 152712 60116
rect 152908 60060 153944 60116
rect 154588 60060 155176 60116
rect 143388 59444 143444 60060
rect 143388 59378 143444 59388
rect 143276 7522 143332 7532
rect 144508 55636 144564 55646
rect 142716 4162 142772 4172
rect 142940 6804 142996 6814
rect 142940 480 142996 6748
rect 144508 5908 144564 55580
rect 144620 11788 144676 60060
rect 146188 59444 146244 59454
rect 146188 56644 146244 59388
rect 146188 56578 146244 56588
rect 146300 56420 146356 60060
rect 147084 59444 147140 60060
rect 147084 59378 147140 59388
rect 146300 56354 146356 56364
rect 144620 11732 144788 11788
rect 144732 8036 144788 11732
rect 144732 7970 144788 7980
rect 147868 5908 147924 60060
rect 144508 5852 144676 5908
rect 136892 476 137256 480
rect 136892 420 136948 476
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 136108 364 136948 420
rect 137004 392 137256 476
rect 137032 -960 137256 392
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 142744 392 142996 480
rect 144620 480 144676 5852
rect 147868 5842 147924 5852
rect 148652 55524 148708 55534
rect 146748 5012 146804 5022
rect 146748 480 146804 4956
rect 148652 5012 148708 55468
rect 149548 6804 149604 60060
rect 151228 59106 151284 59118
rect 151228 59054 151230 59106
rect 151282 59054 151284 59106
rect 151228 55524 151284 59054
rect 151340 55636 151396 60060
rect 152012 59106 152068 60060
rect 152012 59054 152014 59106
rect 152066 59054 152068 59106
rect 152012 59042 152068 59054
rect 151340 55570 151396 55580
rect 151228 55458 151284 55468
rect 149548 6738 149604 6748
rect 152460 7588 152516 7598
rect 148652 4946 148708 4956
rect 150556 4340 150612 4350
rect 148652 4228 148708 4238
rect 148652 480 148708 4172
rect 150556 480 150612 4284
rect 152460 480 152516 7532
rect 152908 4228 152964 60060
rect 152908 4162 152964 4172
rect 154364 5012 154420 5022
rect 154364 480 154420 4956
rect 154588 4340 154644 60060
rect 156268 59442 156324 59454
rect 156268 59390 156270 59442
rect 156322 59390 156324 59442
rect 156268 5012 156324 59390
rect 156380 7588 156436 60088
rect 156940 60060 157640 60116
rect 157948 60060 158872 60116
rect 159628 60060 160104 60116
rect 161336 60060 161476 60116
rect 156940 59442 156996 60060
rect 156940 59390 156942 59442
rect 156994 59390 156996 59442
rect 156940 59378 156996 59390
rect 156380 7522 156436 7532
rect 156268 4946 156324 4956
rect 154588 4274 154644 4284
rect 156156 4900 156212 4910
rect 156156 480 156212 4844
rect 157948 4900 158004 60060
rect 157948 4834 158004 4844
rect 158172 5012 158228 5022
rect 158172 480 158228 4956
rect 159628 5012 159684 60060
rect 161308 59218 161364 59230
rect 161308 59166 161310 59218
rect 161362 59166 161364 59218
rect 159628 4946 159684 4956
rect 160076 5012 160132 5022
rect 160076 480 160132 4956
rect 144620 392 144872 480
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 392
rect 144648 -960 144872 392
rect 146552 392 146804 480
rect 148456 392 148708 480
rect 150360 392 150612 480
rect 152264 392 152516 480
rect 154168 392 154420 480
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157976 392 158228 480
rect 159880 392 160132 480
rect 161308 420 161364 59166
rect 161420 5012 161476 60060
rect 161868 60060 162568 60116
rect 162988 60060 163800 60116
rect 164668 60060 165032 60116
rect 165340 60060 166264 60116
rect 166348 60060 167496 60116
rect 168028 60060 168728 60116
rect 169708 60060 169960 60116
rect 170156 60060 171192 60116
rect 171612 60060 172424 60116
rect 173068 60060 173656 60116
rect 174748 60060 174888 60116
rect 175084 60060 176120 60116
rect 176652 60060 177352 60116
rect 178108 60060 178584 60116
rect 161868 59218 161924 60060
rect 161868 59166 161870 59218
rect 161922 59166 161924 59218
rect 161868 59154 161924 59166
rect 161420 4946 161476 4956
rect 161644 480 161812 532
rect 161644 476 162008 480
rect 161644 420 161700 476
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161308 364 161700 420
rect 161756 392 162008 476
rect 161784 -960 162008 392
rect 162988 420 163044 60060
rect 163548 480 163716 532
rect 163548 476 163912 480
rect 163548 420 163604 476
rect 162988 364 163604 420
rect 163660 392 163912 476
rect 163688 -960 163912 392
rect 164668 420 164724 60060
rect 165340 58828 165396 60060
rect 164780 58772 165396 58828
rect 164780 55524 164836 58772
rect 164780 55458 164836 55468
rect 166348 5012 166404 60060
rect 166348 4946 166404 4956
rect 166460 55524 166516 55534
rect 165452 480 165620 532
rect 165452 476 165816 480
rect 165452 420 165508 476
rect 164668 364 165508 420
rect 165564 392 165816 476
rect 165592 -960 165816 392
rect 166460 420 166516 55468
rect 168028 55524 168084 60060
rect 168028 55458 168084 55468
rect 169372 5012 169428 5022
rect 167356 480 167524 532
rect 169372 480 169428 4956
rect 169708 5012 169764 60060
rect 170156 58828 170212 60060
rect 169708 4946 169764 4956
rect 169932 58772 170212 58828
rect 169932 4900 169988 58772
rect 171612 56420 171668 60060
rect 171612 56354 171668 56364
rect 169932 4834 169988 4844
rect 171388 55524 171444 55534
rect 171388 480 171444 55468
rect 173068 4452 173124 60060
rect 173068 4386 173124 4396
rect 173180 5012 173236 5022
rect 173180 480 173236 4956
rect 174748 4564 174804 60060
rect 175084 58828 175140 60060
rect 174860 58772 175140 58828
rect 174860 56308 174916 58772
rect 174860 56242 174916 56252
rect 176428 56420 176484 56430
rect 174748 4498 174804 4508
rect 175084 4900 175140 4910
rect 175084 480 175140 4844
rect 167356 476 167720 480
rect 167356 420 167412 476
rect 166460 364 167412 420
rect 167468 392 167720 476
rect 169372 392 169624 480
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 176428 420 176484 56364
rect 176652 55524 176708 60060
rect 176652 55458 176708 55468
rect 178108 4228 178164 60060
rect 178892 55524 178948 55534
rect 178892 4900 178948 55468
rect 178892 4834 178948 4844
rect 178108 4162 178164 4172
rect 178892 4452 178948 4462
rect 176876 480 177044 532
rect 178892 480 178948 4396
rect 179788 4340 179844 60088
rect 179900 60060 181048 60116
rect 181468 60060 182280 60116
rect 183148 60060 183512 60116
rect 183820 60060 184744 60116
rect 184828 60060 185976 60116
rect 186508 60060 187208 60116
rect 188188 60060 188440 60116
rect 188636 60060 189672 60116
rect 189868 60060 190904 60116
rect 191548 60060 192136 60116
rect 193368 60060 193508 60116
rect 179900 5908 179956 60060
rect 179900 5842 179956 5852
rect 180572 56308 180628 56318
rect 180572 5012 180628 56252
rect 181468 7588 181524 60060
rect 181468 7522 181524 7532
rect 180572 4946 180628 4956
rect 182700 5012 182756 5022
rect 179788 4274 179844 4284
rect 180796 4564 180852 4574
rect 180796 480 180852 4508
rect 182700 480 182756 4956
rect 183148 5012 183204 60060
rect 183820 58828 183876 60060
rect 183260 58772 183876 58828
rect 183260 55524 183316 58772
rect 184828 56308 184884 60060
rect 184828 56242 184884 56252
rect 183260 55458 183316 55468
rect 185612 55524 185668 55534
rect 185612 6244 185668 55468
rect 185612 6178 185668 6188
rect 183148 4946 183204 4956
rect 184604 4900 184660 4910
rect 184604 480 184660 4844
rect 186508 4564 186564 60060
rect 188188 4900 188244 60060
rect 188636 58828 188692 60060
rect 188412 58772 188692 58828
rect 188412 11788 188468 58772
rect 188412 11732 188580 11788
rect 188188 4834 188244 4844
rect 186508 4498 186564 4508
rect 188524 4452 188580 11732
rect 189868 4676 189924 60060
rect 190652 56308 190708 56318
rect 190652 6356 190708 56252
rect 190652 6290 190708 6300
rect 189868 4610 189924 4620
rect 190316 5908 190372 5918
rect 188524 4386 188580 4396
rect 188412 4340 188468 4350
rect 186508 4228 186564 4238
rect 186508 480 186564 4172
rect 188412 480 188468 4284
rect 190316 480 190372 5852
rect 191548 4340 191604 60060
rect 193228 59444 193284 59454
rect 191548 4274 191604 4284
rect 192220 7588 192276 7598
rect 192220 480 192276 7532
rect 193228 4228 193284 59388
rect 193452 4788 193508 60060
rect 193900 60060 194600 60116
rect 194908 60060 195832 60116
rect 196588 60060 197064 60116
rect 198296 60060 198436 60116
rect 193900 59444 193956 60060
rect 193900 59378 193956 59388
rect 194908 6020 194964 60060
rect 196588 7812 196644 60060
rect 198268 58994 198324 59006
rect 198268 58942 198270 58994
rect 198322 58942 198324 58994
rect 198268 10948 198324 58942
rect 198380 12740 198436 60060
rect 198828 60060 199528 60116
rect 199948 60060 200760 60116
rect 201628 60060 201992 60116
rect 202300 60060 203224 60116
rect 203308 60060 204456 60116
rect 204988 60060 205688 60116
rect 206668 60060 206920 60116
rect 207340 60060 208152 60116
rect 208348 60060 209384 60116
rect 210028 60060 210616 60116
rect 198828 58994 198884 60060
rect 198828 58942 198830 58994
rect 198882 58942 198884 58994
rect 198828 58930 198884 58942
rect 199948 55636 200004 60060
rect 199948 55570 200004 55580
rect 198380 12674 198436 12684
rect 198268 10882 198324 10892
rect 196588 7746 196644 7756
rect 197932 6356 197988 6366
rect 194908 5954 194964 5964
rect 196028 6244 196084 6254
rect 193452 4722 193508 4732
rect 194124 5012 194180 5022
rect 193228 4162 193284 4172
rect 194124 480 194180 4956
rect 196028 480 196084 6188
rect 197932 480 197988 6300
rect 199948 4564 200004 4574
rect 199948 480 200004 4508
rect 201628 4564 201684 60060
rect 202300 58828 202356 60060
rect 201740 58772 202356 58828
rect 201740 55524 201796 58772
rect 203308 56532 203364 60060
rect 203308 56466 203364 56476
rect 201740 55458 201796 55468
rect 202412 55636 202468 55646
rect 202412 14308 202468 55580
rect 202412 14242 202468 14252
rect 204092 55524 204148 55534
rect 204092 7588 204148 55468
rect 204092 7522 204148 7532
rect 201628 4498 201684 4508
rect 201740 4900 201796 4910
rect 201740 480 201796 4844
rect 203644 4452 203700 4462
rect 203644 480 203700 4396
rect 204988 4452 205044 60060
rect 206668 5908 206724 60060
rect 207340 58828 207396 60060
rect 206780 58772 207396 58828
rect 206780 55524 206836 58772
rect 206780 55458 206836 55468
rect 206668 5842 206724 5852
rect 204988 4386 205044 4396
rect 205548 4676 205604 4686
rect 205548 480 205604 4620
rect 207452 4340 207508 4350
rect 207452 480 207508 4284
rect 208348 4340 208404 60060
rect 210028 56420 210084 60060
rect 211708 59442 211764 59454
rect 211708 59390 211710 59442
rect 211762 59390 211764 59442
rect 210028 56354 210084 56364
rect 210812 56532 210868 56542
rect 209132 55524 209188 55534
rect 209132 16212 209188 55468
rect 209132 16146 209188 16156
rect 210812 6132 210868 56476
rect 210812 6066 210868 6076
rect 208348 4274 208404 4284
rect 209356 4788 209412 4798
rect 209356 480 209412 4732
rect 211260 4228 211316 4238
rect 211260 480 211316 4172
rect 211708 4228 211764 59390
rect 211820 56532 211876 60088
rect 212380 60060 213080 60116
rect 213388 60060 214312 60116
rect 215068 60060 215544 60116
rect 212380 59442 212436 60060
rect 212380 59390 212382 59442
rect 212434 59390 212436 59442
rect 212380 59378 212436 59390
rect 211820 56466 211876 56476
rect 213388 56308 213444 60060
rect 213388 56242 213444 56252
rect 214172 56420 214228 56430
rect 214172 7700 214228 56364
rect 215068 12628 215124 60060
rect 215068 12562 215124 12572
rect 215852 12740 215908 12750
rect 214172 7634 214228 7644
rect 215068 7812 215124 7822
rect 211708 4162 211764 4172
rect 213164 6020 213220 6030
rect 213164 480 213220 5964
rect 215068 480 215124 7756
rect 215852 5012 215908 12684
rect 216748 9380 216804 60088
rect 216860 60060 218008 60116
rect 218428 60060 219240 60116
rect 220220 60060 220472 60116
rect 221004 60060 221704 60116
rect 221788 60060 222936 60116
rect 223468 60060 224168 60116
rect 225260 60060 225400 60116
rect 225932 60060 226632 60116
rect 226828 60060 227864 60116
rect 228508 60060 229096 60116
rect 216860 11396 216916 60060
rect 218428 56420 218484 60060
rect 218428 56354 218484 56364
rect 220108 59444 220164 59454
rect 220108 14644 220164 59388
rect 220220 16100 220276 60060
rect 221004 59444 221060 60060
rect 221004 59378 221060 59388
rect 221788 56644 221844 60060
rect 221788 56578 221844 56588
rect 220220 16034 220276 16044
rect 220108 14578 220164 14588
rect 216860 11330 216916 11340
rect 220108 14308 220164 14318
rect 216748 9314 216804 9324
rect 218316 10948 218372 10958
rect 215852 4946 215908 4956
rect 216972 5012 217028 5022
rect 218316 5012 218372 10892
rect 218316 4956 218484 5012
rect 216972 480 217028 4956
rect 176876 476 177240 480
rect 176876 420 176932 476
rect 176428 364 176932 420
rect 176988 392 177240 476
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 205548 392 205800 480
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218428 420 218484 4956
rect 218764 480 218932 532
rect 218764 476 219128 480
rect 218764 420 218820 476
rect 218428 364 218820 420
rect 218876 392 219128 476
rect 218904 -960 219128 392
rect 220108 420 220164 14252
rect 223468 4676 223524 60060
rect 225148 59218 225204 59230
rect 225148 59166 225150 59218
rect 225202 59166 225204 59218
rect 224252 56420 224308 56430
rect 224252 29428 224308 56364
rect 224252 29362 224308 29372
rect 225148 10948 225204 59166
rect 225260 56420 225316 60060
rect 225932 59218 225988 60060
rect 225932 59166 225934 59218
rect 225986 59166 225988 59218
rect 225932 59154 225988 59166
rect 225260 56354 225316 56364
rect 225148 10882 225204 10892
rect 223468 4610 223524 4620
rect 224588 7588 224644 7598
rect 222684 4564 222740 4574
rect 220668 480 220836 532
rect 222684 480 222740 4508
rect 224588 480 224644 7532
rect 226492 6132 226548 6142
rect 226492 480 226548 6076
rect 226828 4564 226884 60060
rect 227612 56644 227668 56654
rect 227612 6020 227668 56588
rect 228508 7588 228564 60060
rect 230188 59442 230244 59454
rect 230188 59390 230190 59442
rect 230242 59390 230244 59442
rect 228508 7522 228564 7532
rect 229292 56532 229348 56542
rect 229292 6132 229348 56476
rect 229292 6066 229348 6076
rect 227612 5954 227668 5964
rect 226828 4498 226884 4508
rect 228508 4452 228564 4462
rect 228508 480 228564 4396
rect 230188 4452 230244 59390
rect 230300 26068 230356 60088
rect 230860 60060 231560 60116
rect 231868 60060 232792 60116
rect 233548 60060 234024 60116
rect 230860 59442 230916 60060
rect 230860 59390 230862 59442
rect 230914 59390 230916 59442
rect 230860 59378 230916 59390
rect 230300 26002 230356 26012
rect 231868 15988 231924 60060
rect 231868 15922 231924 15932
rect 231980 16212 232036 16222
rect 231980 11788 232036 16156
rect 231980 11732 232260 11788
rect 230188 4386 230244 4396
rect 230300 5908 230356 5918
rect 230300 480 230356 5852
rect 232204 480 232260 11732
rect 233548 5908 233604 60060
rect 234332 56308 234388 56318
rect 234332 6244 234388 56252
rect 235228 9268 235284 60088
rect 235340 60060 236488 60116
rect 236908 60060 237720 60116
rect 238700 60060 238952 60116
rect 239484 60060 240184 60116
rect 240268 60060 241416 60116
rect 241948 60060 242648 60116
rect 243628 60060 243880 60116
rect 244300 60060 245112 60116
rect 245308 60060 246344 60116
rect 246988 60060 247576 60116
rect 248668 60060 248808 60116
rect 249004 60060 250040 60116
rect 250348 60060 251272 60116
rect 252028 60060 252504 60116
rect 235340 56308 235396 60060
rect 236908 56756 236964 60060
rect 236908 56690 236964 56700
rect 238588 59444 238644 59454
rect 235340 56242 235396 56252
rect 238588 12740 238644 59388
rect 238700 47908 238756 60060
rect 239484 59444 239540 60060
rect 239484 59378 239540 59388
rect 240268 55524 240324 60060
rect 240268 55458 240324 55468
rect 238700 47842 238756 47852
rect 241948 18004 242004 60060
rect 241948 17938 242004 17948
rect 242732 56756 242788 56766
rect 242732 17668 242788 56700
rect 242732 17602 242788 17612
rect 238588 12674 238644 12684
rect 235228 9202 235284 9212
rect 234332 6178 234388 6188
rect 236012 7700 236068 7710
rect 233548 5842 233604 5852
rect 234108 4340 234164 4350
rect 234108 480 234164 4284
rect 236012 480 236068 7644
rect 243628 7700 243684 60060
rect 244300 58828 244356 60060
rect 243740 58772 244356 58828
rect 243740 36148 243796 58772
rect 243740 36082 243796 36092
rect 243628 7634 243684 7644
rect 243740 12628 243796 12638
rect 241724 6244 241780 6254
rect 237916 6132 237972 6142
rect 237916 480 237972 6076
rect 239820 4228 239876 4238
rect 239820 480 239876 4172
rect 241724 480 241780 6188
rect 243740 480 243796 12572
rect 245308 4340 245364 60060
rect 246092 55524 246148 55534
rect 246092 21028 246148 55468
rect 246092 20962 246148 20972
rect 246988 11172 247044 60060
rect 246988 11106 247044 11116
rect 247436 11396 247492 11406
rect 245308 4274 245364 4284
rect 245532 9380 245588 9390
rect 245532 480 245588 9324
rect 247436 480 247492 11340
rect 248668 2548 248724 60060
rect 249004 58828 249060 60060
rect 248780 58772 249060 58828
rect 248780 56532 248836 58772
rect 248780 56466 248836 56476
rect 248668 2482 248724 2492
rect 248780 29428 248836 29438
rect 220668 476 221032 480
rect 220668 420 220724 476
rect 220108 364 220724 420
rect 220780 392 221032 476
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 234108 392 234360 480
rect 236012 392 236264 480
rect 237916 392 238168 480
rect 239820 392 240072 480
rect 241724 392 241976 480
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 392
rect 243656 -960 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 248780 420 248836 29372
rect 250348 19348 250404 60060
rect 250348 19282 250404 19292
rect 251132 56420 251188 56430
rect 250348 16100 250404 16110
rect 249228 480 249396 532
rect 249228 476 249592 480
rect 249228 420 249284 476
rect 248780 364 249284 420
rect 249340 392 249592 476
rect 249368 -960 249592 392
rect 250348 420 250404 16044
rect 251132 6132 251188 56364
rect 252028 14420 252084 60060
rect 252028 14354 252084 14364
rect 252140 14644 252196 14654
rect 251132 6066 251188 6076
rect 251132 480 251300 532
rect 251132 476 251496 480
rect 251132 420 251188 476
rect 250348 364 251188 420
rect 251244 392 251496 476
rect 251272 -960 251496 392
rect 252140 420 252196 14588
rect 253708 4228 253764 60088
rect 253820 60060 254968 60116
rect 255388 60060 256200 60116
rect 257068 60060 257432 60116
rect 257628 60060 258664 60116
rect 258748 60060 259896 60116
rect 260428 60060 261128 60116
rect 262220 60060 262360 60116
rect 262892 60060 263592 60116
rect 263788 60060 264824 60116
rect 265468 60060 266056 60116
rect 267148 60060 267288 60116
rect 267484 60060 268520 60116
rect 268828 60060 269752 60116
rect 270508 60060 270984 60116
rect 253820 56420 253876 60060
rect 255388 56756 255444 60060
rect 255388 56690 255444 56700
rect 253820 56354 253876 56364
rect 253708 4162 253764 4172
rect 255052 6020 255108 6030
rect 253036 480 253204 532
rect 255052 480 255108 5964
rect 257068 4900 257124 60060
rect 257628 58828 257684 60060
rect 257180 58772 257684 58828
rect 257180 24388 257236 58772
rect 258748 56868 258804 60060
rect 258748 56802 258804 56812
rect 257180 24322 257236 24332
rect 260428 6244 260484 60060
rect 262108 59218 262164 59230
rect 262108 59166 262110 59218
rect 262162 59166 262164 59218
rect 261212 56756 261268 56766
rect 261212 34468 261268 56700
rect 261212 34402 261268 34412
rect 260428 6178 260484 6188
rect 260764 10948 260820 10958
rect 257068 4834 257124 4844
rect 258860 6132 258916 6142
rect 257068 4676 257124 4686
rect 257068 480 257124 4620
rect 258860 480 258916 6076
rect 260764 480 260820 10892
rect 262108 6132 262164 59166
rect 262220 14308 262276 60060
rect 262892 59218 262948 60060
rect 262892 59166 262894 59218
rect 262946 59166 262948 59218
rect 262892 59154 262948 59166
rect 262220 14242 262276 14252
rect 262108 6066 262164 6076
rect 263788 4788 263844 60060
rect 264572 56868 264628 56878
rect 264572 37828 264628 56812
rect 265468 44548 265524 60060
rect 265468 44482 265524 44492
rect 266252 56532 266308 56542
rect 264572 37762 264628 37772
rect 265468 26068 265524 26078
rect 263788 4722 263844 4732
rect 264572 7588 264628 7598
rect 262668 4564 262724 4574
rect 262668 480 262724 4508
rect 264572 480 264628 7532
rect 253036 476 253400 480
rect 253036 420 253092 476
rect 252140 364 253092 420
rect 253148 392 253400 476
rect 255052 392 255304 480
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 265468 420 265524 26012
rect 266252 7812 266308 56476
rect 267148 16100 267204 60060
rect 267484 58828 267540 60060
rect 267260 58772 267540 58828
rect 267260 56532 267316 58772
rect 267260 56466 267316 56476
rect 267148 16034 267204 16044
rect 267932 56308 267988 56318
rect 266252 7746 266308 7756
rect 267932 6020 267988 56252
rect 268828 12628 268884 60060
rect 268828 12562 268884 12572
rect 268940 15988 268996 15998
rect 267932 5954 267988 5964
rect 268380 4452 268436 4462
rect 266364 480 266532 532
rect 268380 480 268436 4396
rect 266364 476 266728 480
rect 266364 420 266420 476
rect 265468 364 266420 420
rect 266476 392 266728 476
rect 268380 392 268632 480
rect 266504 -960 266728 392
rect 268408 -960 268632 392
rect 268940 420 268996 15932
rect 270508 11060 270564 60060
rect 272188 11788 272244 60088
rect 272300 60060 273448 60116
rect 273868 60060 274680 60116
rect 275548 60060 275912 60116
rect 276220 60060 277144 60116
rect 277228 60060 278376 60116
rect 278908 60060 279608 60116
rect 280588 60060 280840 60116
rect 281260 60060 282072 60116
rect 282268 60060 283304 60116
rect 283948 60060 284536 60116
rect 285628 60060 285768 60116
rect 285964 60060 287000 60116
rect 287308 60060 288232 60116
rect 289100 60060 289464 60116
rect 290696 60060 290948 60116
rect 272300 55524 272356 60060
rect 272300 55458 272356 55468
rect 273868 12852 273924 60060
rect 274652 55524 274708 55534
rect 274652 32788 274708 55468
rect 274652 32722 274708 32732
rect 273868 12786 273924 12796
rect 272188 11732 272356 11788
rect 270508 10994 270564 11004
rect 272188 5908 272244 5918
rect 270172 480 270340 532
rect 272188 480 272244 5852
rect 272300 4676 272356 11732
rect 272300 4610 272356 4620
rect 274092 9268 274148 9278
rect 274092 480 274148 9212
rect 275548 4564 275604 60060
rect 276220 58828 276276 60060
rect 275660 58772 276276 58828
rect 275660 56308 275716 58772
rect 275660 56242 275716 56252
rect 277228 29540 277284 60060
rect 278908 54740 278964 60060
rect 278908 54674 278964 54684
rect 279692 56532 279748 56542
rect 277228 29474 277284 29484
rect 278908 47908 278964 47918
rect 277228 17668 277284 17678
rect 275548 4498 275604 4508
rect 275996 6020 276052 6030
rect 275996 480 276052 5964
rect 270172 476 270536 480
rect 270172 420 270228 476
rect 268940 364 270228 420
rect 270284 392 270536 476
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277228 420 277284 17612
rect 277788 480 277956 532
rect 277788 476 278152 480
rect 277788 420 277844 476
rect 277228 364 277844 420
rect 277900 392 278152 476
rect 277928 -960 278152 392
rect 278908 420 278964 47852
rect 279692 9268 279748 56476
rect 279692 9202 279748 9212
rect 280588 6020 280644 60060
rect 281260 58828 281316 60060
rect 280700 58772 281316 58828
rect 280700 29428 280756 58772
rect 280700 29362 280756 29372
rect 280588 5954 280644 5964
rect 280700 12740 280756 12750
rect 279692 480 279860 532
rect 279692 476 280056 480
rect 279692 420 279748 476
rect 278908 364 279748 420
rect 279804 392 280056 476
rect 279832 -960 280056 392
rect 280700 420 280756 12684
rect 282268 4452 282324 60060
rect 282268 4386 282324 4396
rect 282380 21028 282436 21038
rect 281596 480 281764 532
rect 281596 476 281960 480
rect 281596 420 281652 476
rect 280700 364 281652 420
rect 281708 392 281960 476
rect 281736 -960 281960 392
rect 282380 420 282436 20972
rect 283948 7588 284004 60060
rect 285628 17780 285684 60060
rect 285964 58828 286020 60060
rect 285740 58772 286020 58828
rect 285740 56756 285796 58772
rect 285740 56690 285796 56700
rect 286412 56420 286468 56430
rect 285628 17714 285684 17724
rect 285740 18004 285796 18014
rect 283948 7522 284004 7532
rect 283500 480 283668 532
rect 285740 480 285796 17948
rect 286412 7924 286468 56364
rect 287308 10948 287364 60060
rect 287308 10882 287364 10892
rect 288988 36148 289044 36158
rect 286412 7858 286468 7868
rect 283500 476 283864 480
rect 283500 420 283556 476
rect 282380 364 283556 420
rect 283612 392 283864 476
rect 283640 -960 283864 392
rect 285544 392 285796 480
rect 287420 7700 287476 7710
rect 287420 480 287476 7644
rect 287420 392 287672 480
rect 285544 -960 285768 392
rect 287448 -960 287672 392
rect 288988 420 289044 36092
rect 289100 26180 289156 60060
rect 290668 59332 290724 59342
rect 290668 56532 290724 59276
rect 290892 56644 290948 60060
rect 291228 60060 291928 60116
rect 292348 60060 293160 60116
rect 294252 60060 294392 60116
rect 294924 60060 295624 60116
rect 295708 60060 296856 60116
rect 297388 60060 298088 60116
rect 299180 60060 299320 60116
rect 299852 60060 300552 60116
rect 300748 60060 301784 60116
rect 302428 60060 303016 60116
rect 291228 59332 291284 60060
rect 291228 59266 291284 59276
rect 290892 56578 290948 56588
rect 290668 56466 290724 56476
rect 289100 26114 289156 26124
rect 292348 5908 292404 60060
rect 294028 59444 294084 59454
rect 294028 56420 294084 59388
rect 294028 56354 294084 56364
rect 294252 55524 294308 60060
rect 294924 59444 294980 60060
rect 294924 59378 294980 59388
rect 294252 55458 294308 55468
rect 295708 17668 295764 60060
rect 296492 56644 296548 56654
rect 296492 27860 296548 56588
rect 296492 27794 296548 27804
rect 297388 19572 297444 60060
rect 299068 59218 299124 59230
rect 299068 59166 299070 59218
rect 299122 59166 299124 59218
rect 298172 55524 298228 55534
rect 298172 31220 298228 55468
rect 298172 31154 298228 31164
rect 297388 19506 297444 19516
rect 295708 17602 295764 17612
rect 297388 19348 297444 19358
rect 292348 5842 292404 5852
rect 293132 11172 293188 11182
rect 291228 4340 291284 4350
rect 289212 480 289380 532
rect 291228 480 291284 4284
rect 293132 480 293188 11116
rect 296940 7812 296996 7822
rect 295036 2548 295092 2558
rect 295036 480 295092 2492
rect 296940 480 296996 7756
rect 289212 476 289576 480
rect 289212 420 289268 476
rect 288988 364 289268 420
rect 289324 392 289576 476
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 297388 420 297444 19292
rect 299068 12740 299124 59166
rect 299180 46228 299236 60060
rect 299852 59218 299908 60060
rect 299852 59166 299854 59218
rect 299906 59166 299908 59218
rect 299852 59154 299908 59166
rect 299180 46162 299236 46172
rect 299068 12674 299124 12684
rect 300748 4340 300804 60060
rect 300748 4274 300804 4284
rect 300860 14420 300916 14430
rect 298732 480 298900 532
rect 300860 480 300916 14364
rect 302428 7812 302484 60060
rect 302428 7746 302484 7756
rect 304108 59108 304164 59118
rect 302652 4228 302708 4238
rect 302652 480 302708 4172
rect 304108 4228 304164 59052
rect 304220 26068 304276 60088
rect 304780 60060 305480 60116
rect 305788 60060 306712 60116
rect 307468 60060 307944 60116
rect 304780 59108 304836 60060
rect 304780 59042 304836 59052
rect 304220 26002 304276 26012
rect 305788 15988 305844 60060
rect 305788 15922 305844 15932
rect 305900 34468 305956 34478
rect 304108 4162 304164 4172
rect 304556 7924 304612 7934
rect 304556 480 304612 7868
rect 298732 476 299096 480
rect 298732 420 298788 476
rect 297388 364 298788 420
rect 298844 392 299096 476
rect 298872 -960 299096 392
rect 300776 -960 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 305900 420 305956 34412
rect 307468 24612 307524 60060
rect 309148 55524 309204 60088
rect 309372 60060 310408 60116
rect 310828 60060 311640 60116
rect 312620 60060 312872 60116
rect 313404 60060 314104 60116
rect 314188 60060 315336 60116
rect 315868 60060 316568 60116
rect 317660 60060 317800 60116
rect 318332 60060 319032 60116
rect 319228 60060 320264 60116
rect 321132 60060 321496 60116
rect 309372 55860 309428 60060
rect 309372 55794 309428 55804
rect 309148 55458 309204 55468
rect 310828 48020 310884 60060
rect 312508 59444 312564 59454
rect 310828 47954 310884 47964
rect 311612 55524 311668 55534
rect 307468 24546 307524 24556
rect 310828 37828 310884 37838
rect 308252 24388 308308 24398
rect 308252 5012 308308 24332
rect 308252 4946 308308 4956
rect 310268 5012 310324 5022
rect 308364 4900 308420 4910
rect 306348 480 306516 532
rect 308364 480 308420 4844
rect 310268 480 310324 4956
rect 306348 476 306712 480
rect 306348 420 306404 476
rect 305900 364 306404 420
rect 306460 392 306712 476
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 310828 420 310884 37772
rect 311612 37828 311668 55468
rect 312508 54628 312564 59388
rect 312620 55524 312676 60060
rect 313404 59444 313460 60060
rect 313404 59378 313460 59388
rect 312620 55458 312676 55468
rect 312508 54562 312564 54572
rect 311612 37762 311668 37772
rect 314188 19348 314244 60060
rect 314972 55524 315028 55534
rect 314972 36148 315028 55468
rect 314972 36082 315028 36092
rect 314188 19282 314244 19292
rect 315868 14644 315924 60060
rect 317548 59218 317604 59230
rect 317548 59166 317550 59218
rect 317602 59166 317604 59218
rect 315980 55860 316036 55870
rect 315980 49588 316036 55804
rect 315980 49522 316036 49532
rect 317548 27748 317604 59166
rect 317660 56644 317716 60060
rect 318332 59218 318388 60060
rect 318332 59166 318334 59218
rect 318386 59166 318388 59218
rect 318332 59154 318388 59166
rect 317660 56578 317716 56588
rect 317548 27682 317604 27692
rect 315868 14578 315924 14588
rect 315868 14308 315924 14318
rect 315868 11788 315924 14252
rect 315868 11732 316036 11788
rect 314188 6244 314244 6254
rect 312060 480 312228 532
rect 314188 480 314244 6188
rect 315980 480 316036 11732
rect 319228 11172 319284 60060
rect 319228 11106 319284 11116
rect 320908 44548 320964 44558
rect 317884 6132 317940 6142
rect 317884 480 317940 6076
rect 319788 4788 319844 4798
rect 319788 480 319844 4732
rect 312060 476 312424 480
rect 312060 420 312116 476
rect 310828 364 312116 420
rect 312172 392 312424 476
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 320908 420 320964 44492
rect 321132 44548 321188 60060
rect 321132 44482 321188 44492
rect 322588 59442 322644 59454
rect 322588 59390 322590 59442
rect 322642 59390 322644 59442
rect 322588 14308 322644 59390
rect 322700 31108 322756 60088
rect 323260 60060 323960 60116
rect 324268 60060 325192 60116
rect 325948 60060 326424 60116
rect 323260 59442 323316 60060
rect 323260 59390 323262 59442
rect 323314 59390 323316 59442
rect 323260 59378 323316 59390
rect 322700 31042 322756 31052
rect 322588 14242 322644 14252
rect 322700 16100 322756 16110
rect 321580 480 321748 532
rect 321580 476 321944 480
rect 321580 420 321636 476
rect 320908 364 321636 420
rect 321692 392 321944 476
rect 321720 -960 321944 392
rect 322700 420 322756 16044
rect 324268 7700 324324 60060
rect 325052 56756 325108 56766
rect 325052 18004 325108 56700
rect 325948 56756 326004 60060
rect 325948 56690 326004 56700
rect 325052 17938 325108 17948
rect 325948 12628 326004 12638
rect 324268 7634 324324 7644
rect 325500 9268 325556 9278
rect 323484 480 323652 532
rect 325500 480 325556 9212
rect 323484 476 323848 480
rect 323484 420 323540 476
rect 322700 364 323540 420
rect 323596 392 323848 476
rect 325500 392 325752 480
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 325948 420 326004 12572
rect 327628 12628 327684 60088
rect 327740 60060 328888 60116
rect 329308 60060 330120 60116
rect 330988 60060 331352 60116
rect 331884 60060 332584 60116
rect 332668 60060 333816 60116
rect 334348 60060 335048 60116
rect 336140 60060 336280 60116
rect 336812 60060 337512 60116
rect 337708 60060 338744 60116
rect 339388 60060 339976 60116
rect 327740 32900 327796 60060
rect 327740 32834 327796 32844
rect 327628 12562 327684 12572
rect 329308 11788 329364 60060
rect 330092 56756 330148 56766
rect 329308 11732 329476 11788
rect 329308 11060 329364 11070
rect 327292 480 327460 532
rect 329308 480 329364 11004
rect 329420 6244 329476 11732
rect 330092 9380 330148 56700
rect 330988 55524 331044 60060
rect 331884 58828 331940 60060
rect 331212 58772 331940 58828
rect 331212 56756 331268 58772
rect 331212 56690 331268 56700
rect 330988 55458 331044 55468
rect 332668 22820 332724 60060
rect 333452 55524 333508 55534
rect 333452 38052 333508 55468
rect 334348 39508 334404 60060
rect 336028 59218 336084 59230
rect 336028 59166 336030 59218
rect 336082 59166 336084 59218
rect 334348 39442 334404 39452
rect 335132 56308 335188 56318
rect 333452 37986 333508 37996
rect 332668 22754 332724 22764
rect 332780 32788 332836 32798
rect 330092 9314 330148 9324
rect 329420 6178 329476 6188
rect 331212 4676 331268 4686
rect 331212 480 331268 4620
rect 327292 476 327656 480
rect 327292 420 327348 476
rect 325948 364 327348 420
rect 327404 392 327656 476
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 332780 420 332836 32732
rect 334348 12852 334404 12862
rect 333004 480 333172 532
rect 333004 476 333368 480
rect 333004 420 333060 476
rect 332780 364 333060 420
rect 333116 392 333368 476
rect 333144 -960 333368 392
rect 334348 420 334404 12796
rect 335132 5796 335188 56252
rect 336028 11060 336084 59166
rect 336140 56308 336196 60060
rect 336812 59218 336868 60060
rect 336812 59166 336814 59218
rect 336866 59166 336868 59218
rect 336812 59154 336868 59166
rect 336140 56242 336196 56252
rect 337708 12852 337764 60060
rect 337708 12786 337764 12796
rect 336028 10994 336084 11004
rect 335132 5730 335188 5740
rect 338828 5796 338884 5806
rect 336924 4564 336980 4574
rect 334908 480 335076 532
rect 336924 480 336980 4508
rect 338828 480 338884 5740
rect 339388 2660 339444 60060
rect 341068 59444 341124 59454
rect 339388 2594 339444 2604
rect 339500 29540 339556 29550
rect 334908 476 335272 480
rect 334908 420 334964 476
rect 334348 364 334964 420
rect 335020 392 335272 476
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 339500 420 339556 29484
rect 341068 6132 341124 59388
rect 341180 21140 341236 60088
rect 341740 60060 342440 60116
rect 342860 60060 343672 60116
rect 344428 60060 344904 60116
rect 341740 59444 341796 60060
rect 341740 59378 341796 59388
rect 341180 21074 341236 21084
rect 342748 54740 342804 54750
rect 341068 6066 341124 6076
rect 340620 480 340788 532
rect 342748 480 342804 54684
rect 342860 46452 342916 60060
rect 344428 56868 344484 60060
rect 344428 56802 344484 56812
rect 342860 46386 342916 46396
rect 346108 34580 346164 60088
rect 346220 60060 347368 60116
rect 347788 60060 348600 60116
rect 349580 60060 349832 60116
rect 350364 60060 351064 60116
rect 351148 60060 352296 60116
rect 352828 60060 353528 60116
rect 354620 60060 354760 60116
rect 355292 60060 355992 60116
rect 356188 60060 357224 60116
rect 357868 60060 358456 60116
rect 346220 44772 346276 60060
rect 347788 54964 347844 60060
rect 347788 54898 347844 54908
rect 349468 59444 349524 59454
rect 346220 44706 346276 44716
rect 346108 34514 346164 34524
rect 346108 29428 346164 29438
rect 344540 6020 344596 6030
rect 344540 480 344596 5964
rect 340620 476 340984 480
rect 340620 420 340676 476
rect 339500 364 340676 420
rect 340732 392 340984 476
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 344568 -960 344792 392
rect 346108 420 346164 29372
rect 349468 16100 349524 59388
rect 349580 53172 349636 60060
rect 350364 59444 350420 60060
rect 350364 59378 350420 59388
rect 349580 53106 349636 53116
rect 351148 29540 351204 60060
rect 351148 29474 351204 29484
rect 351932 56756 351988 56766
rect 351932 17892 351988 56700
rect 352828 19460 352884 60060
rect 354508 59218 354564 59230
rect 354508 59166 354510 59218
rect 354562 59166 354564 59218
rect 354508 36260 354564 59166
rect 354620 58100 354676 60060
rect 355292 59218 355348 60060
rect 355292 59166 355294 59218
rect 355346 59166 355348 59218
rect 355292 59154 355348 59166
rect 354620 58034 354676 58044
rect 354508 36194 354564 36204
rect 355292 56868 355348 56878
rect 352828 19394 352884 19404
rect 351932 17826 351988 17836
rect 352828 18004 352884 18014
rect 349468 16034 349524 16044
rect 351148 17780 351204 17790
rect 350252 7588 350308 7598
rect 348348 4452 348404 4462
rect 346332 480 346500 532
rect 348348 480 348404 4396
rect 350252 480 350308 7532
rect 346332 476 346696 480
rect 346332 420 346388 476
rect 346108 364 346388 420
rect 346444 392 346696 476
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 351148 420 351204 17724
rect 352044 480 352212 532
rect 352044 476 352408 480
rect 352044 420 352100 476
rect 351148 364 352100 420
rect 352156 392 352408 476
rect 352184 -960 352408 392
rect 352828 420 352884 17948
rect 355292 17780 355348 56812
rect 356188 48132 356244 60060
rect 356188 48066 356244 48076
rect 356972 56532 357028 56542
rect 355292 17714 355348 17724
rect 355964 10948 356020 10958
rect 353948 480 354116 532
rect 355964 480 356020 10892
rect 356972 8148 357028 56476
rect 357868 41412 357924 60060
rect 357868 41346 357924 41356
rect 359548 59442 359604 59454
rect 359548 59390 359550 59442
rect 359602 59390 359604 59442
rect 359548 39620 359604 59390
rect 359660 51492 359716 60088
rect 360220 60060 360920 60116
rect 361228 60060 362152 60116
rect 362908 60060 363384 60116
rect 360220 59442 360276 60060
rect 360220 59390 360222 59442
rect 360274 59390 360276 59442
rect 360220 59378 360276 59390
rect 359660 51426 359716 51436
rect 359548 39554 359604 39564
rect 359548 27860 359604 27870
rect 356972 8082 357028 8092
rect 357868 26180 357924 26190
rect 357868 480 357924 26124
rect 359548 11788 359604 27804
rect 361228 21028 361284 60060
rect 361228 20962 361284 20972
rect 362012 56420 362068 56430
rect 359548 11732 359828 11788
rect 359772 480 359828 11732
rect 361676 8148 361732 8158
rect 361676 480 361732 8092
rect 362012 6356 362068 56364
rect 362908 56420 362964 60060
rect 362908 56354 362964 56364
rect 362012 6290 362068 6300
rect 364588 6020 364644 60088
rect 364700 60060 365848 60116
rect 366268 60060 367080 60116
rect 367948 60060 368312 60116
rect 368620 60060 369544 60116
rect 369628 60060 370776 60116
rect 371308 60060 372008 60116
rect 373100 60060 373240 60116
rect 373772 60060 374472 60116
rect 374668 60060 375704 60116
rect 376348 60060 376936 60116
rect 364700 56532 364756 60060
rect 366268 56868 366324 60060
rect 366268 56802 366324 56812
rect 364700 56466 364756 56476
rect 365596 56420 365652 56430
rect 365596 51380 365652 56364
rect 365596 51314 365652 51324
rect 364588 5954 364644 5964
rect 364700 31220 364756 31230
rect 363580 5908 363636 5918
rect 363580 480 363636 5852
rect 353948 476 354312 480
rect 353948 420 354004 476
rect 352828 364 354004 420
rect 354060 392 354312 476
rect 355964 392 356216 480
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 363580 392 363832 480
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 -960 363832 392
rect 364700 420 364756 31164
rect 367948 26180 368004 60060
rect 368620 58828 368676 60060
rect 368060 58772 368676 58828
rect 368060 46340 368116 58772
rect 368060 46274 368116 46284
rect 369628 29428 369684 60060
rect 369628 29362 369684 29372
rect 370412 56644 370468 56654
rect 367948 26114 368004 26124
rect 367948 17668 368004 17678
rect 367388 6356 367444 6366
rect 365372 480 365540 532
rect 367388 480 367444 6300
rect 365372 476 365736 480
rect 365372 420 365428 476
rect 364700 364 365428 420
rect 365484 392 365736 476
rect 367388 392 367640 480
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 367948 420 368004 17612
rect 370412 7924 370468 56588
rect 371308 31220 371364 60060
rect 372988 59218 373044 59230
rect 372988 59166 372990 59218
rect 373042 59166 373044 59218
rect 372092 56868 372148 56878
rect 372092 42980 372148 56812
rect 372092 42914 372148 42924
rect 371308 31154 371364 31164
rect 370412 7858 370468 7868
rect 371308 19572 371364 19582
rect 369180 480 369348 532
rect 371308 480 371364 19516
rect 372988 7588 373044 59166
rect 373100 53060 373156 60060
rect 373772 59218 373828 60060
rect 373772 59166 373774 59218
rect 373826 59166 373828 59218
rect 373772 59154 373828 59166
rect 373100 52994 373156 53004
rect 374668 34468 374724 60060
rect 374668 34402 374724 34412
rect 374780 46228 374836 46238
rect 372988 7522 373044 7532
rect 374668 12740 374724 12750
rect 373324 5012 373380 5022
rect 373324 480 373380 4956
rect 369180 476 369544 480
rect 369180 420 369236 476
rect 367948 364 369236 420
rect 369292 392 369544 476
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373128 392 373380 480
rect 374668 420 374724 12684
rect 374780 5012 374836 46172
rect 374780 4946 374836 4956
rect 376348 2548 376404 60060
rect 378028 59442 378084 59454
rect 378028 59390 378030 59442
rect 378082 59390 378084 59442
rect 378028 9268 378084 59390
rect 378140 57988 378196 60088
rect 378700 60060 379400 60116
rect 379708 60060 380632 60116
rect 381388 60060 381864 60116
rect 383096 60060 383236 60116
rect 378700 59442 378756 60060
rect 378700 59390 378702 59442
rect 378754 59390 378756 59442
rect 378700 59378 378756 59390
rect 378140 57922 378196 57932
rect 379708 22708 379764 60060
rect 381388 55524 381444 60060
rect 381388 55458 381444 55468
rect 383068 59218 383124 59230
rect 383068 59166 383070 59218
rect 383122 59166 383124 59218
rect 379708 22642 379764 22652
rect 379820 26068 379876 26078
rect 378028 9202 378084 9212
rect 378812 7812 378868 7822
rect 376348 2482 376404 2492
rect 376908 4340 376964 4350
rect 374892 480 375060 532
rect 376908 480 376964 4284
rect 378812 480 378868 7756
rect 374892 476 375256 480
rect 374892 420 374948 476
rect 373128 -960 373352 392
rect 374668 364 374948 420
rect 375004 392 375256 476
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 379820 420 379876 26012
rect 383068 24500 383124 59166
rect 383180 56644 383236 60060
rect 383628 60060 384328 60116
rect 384748 60060 385560 60116
rect 386540 60060 386792 60116
rect 387324 60060 388024 60116
rect 388332 60060 389256 60116
rect 389900 60060 390488 60116
rect 391580 60060 391720 60116
rect 392252 60060 392952 60116
rect 393148 60060 394184 60116
rect 394940 60060 395416 60116
rect 383628 59218 383684 60060
rect 383628 59166 383630 59218
rect 383682 59166 383684 59218
rect 383628 59154 383684 59166
rect 384748 56756 384804 60060
rect 384748 56690 384804 56700
rect 386428 59444 386484 59454
rect 383180 56578 383236 56588
rect 383852 55524 383908 55534
rect 383852 46228 383908 55468
rect 383852 46162 383908 46172
rect 383068 24434 383124 24444
rect 386428 24388 386484 59388
rect 386540 56420 386596 60060
rect 387324 59444 387380 60060
rect 387324 59378 387380 59388
rect 386540 56354 386596 56364
rect 388332 37940 388388 60060
rect 388332 37874 388388 37884
rect 389788 49588 389844 49598
rect 388108 37828 388164 37838
rect 386428 24322 386484 24332
rect 386540 24612 386596 24622
rect 383068 15988 383124 15998
rect 382620 4228 382676 4238
rect 380604 480 380772 532
rect 382620 480 382676 4172
rect 380604 476 380968 480
rect 380604 420 380660 476
rect 379820 364 380660 420
rect 380716 392 380968 476
rect 382620 392 382872 480
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 383068 420 383124 15932
rect 384412 480 384580 532
rect 386540 480 386596 24556
rect 388108 11788 388164 37772
rect 388108 11732 388388 11788
rect 388332 480 388388 11732
rect 384412 476 384776 480
rect 384412 420 384468 476
rect 383068 364 384468 420
rect 384524 392 384776 476
rect 384552 -960 384776 392
rect 386456 -960 386680 480
rect 388332 392 388584 480
rect 388360 -960 388584 392
rect 389788 420 389844 49532
rect 389900 47908 389956 60060
rect 391468 59218 391524 59230
rect 391468 59166 391470 59218
rect 391522 59166 391524 59218
rect 390348 56756 390404 56766
rect 390348 49700 390404 56700
rect 390348 49634 390404 49644
rect 389900 47842 389956 47852
rect 391468 10948 391524 59166
rect 391580 55524 391636 60060
rect 392252 59218 392308 60060
rect 392252 59166 392254 59218
rect 392306 59166 392308 59218
rect 392252 59154 392308 59166
rect 393148 56756 393204 60060
rect 393148 56690 393204 56700
rect 391580 55458 391636 55468
rect 393596 56644 393652 56654
rect 391468 10882 391524 10892
rect 391580 48020 391636 48030
rect 390124 480 390292 532
rect 390124 476 390488 480
rect 390124 420 390180 476
rect 389788 364 390180 420
rect 390236 392 390488 476
rect 390264 -960 390488 392
rect 391580 420 391636 47964
rect 393596 48020 393652 56588
rect 393596 47954 393652 47964
rect 393932 55524 393988 55534
rect 393932 44660 393988 55468
rect 393932 44594 393988 44604
rect 394828 54628 394884 54638
rect 393148 36148 393204 36158
rect 392028 480 392196 532
rect 392028 476 392392 480
rect 392028 420 392084 476
rect 391580 364 392084 420
rect 392140 392 392392 476
rect 392168 -960 392392 392
rect 393148 420 393204 36092
rect 393932 480 394100 532
rect 393932 476 394296 480
rect 393932 420 393988 476
rect 393148 364 393988 420
rect 394044 392 394296 476
rect 394072 -960 394296 392
rect 394828 420 394884 54572
rect 394940 32788 394996 60060
rect 394940 32722 394996 32732
rect 396508 59442 396564 59454
rect 396508 59390 396510 59442
rect 396562 59390 396564 59442
rect 396508 17668 396564 59390
rect 396620 51268 396676 60088
rect 397180 60060 397880 60116
rect 398188 60060 399112 60116
rect 399868 60060 400344 60116
rect 401576 60060 401716 60116
rect 397180 59442 397236 60060
rect 397180 59390 397182 59442
rect 397234 59390 397236 59442
rect 397180 59378 397236 59390
rect 398188 56644 398244 60060
rect 398188 56578 398244 56588
rect 396620 51202 396676 51212
rect 396508 17602 396564 17612
rect 396620 19348 396676 19358
rect 395836 480 396004 532
rect 395836 476 396200 480
rect 395836 420 395892 476
rect 394828 364 395892 420
rect 395948 392 396200 476
rect 395976 -960 396200 392
rect 396620 420 396676 19292
rect 399868 14420 399924 60060
rect 401548 59218 401604 59230
rect 401548 59166 401550 59218
rect 401602 59166 401604 59218
rect 401548 37828 401604 59166
rect 401660 55524 401716 60060
rect 402108 60060 402808 60116
rect 403228 60060 404040 60116
rect 404908 60060 405272 60116
rect 405468 60060 406504 60116
rect 406700 60060 407736 60116
rect 408268 60060 408968 60116
rect 410060 60060 410200 60116
rect 410732 60060 411432 60116
rect 411628 60060 412664 60116
rect 413308 60060 413896 60116
rect 402108 59218 402164 60060
rect 402108 59166 402110 59218
rect 402162 59166 402164 59218
rect 402108 59154 402164 59166
rect 401660 55458 401716 55468
rect 403228 49588 403284 60060
rect 403228 49522 403284 49532
rect 401548 37762 401604 37772
rect 403228 27748 403284 27758
rect 399868 14354 399924 14364
rect 399980 14644 400036 14654
rect 397740 480 397908 532
rect 399980 480 400036 14588
rect 397740 476 398104 480
rect 397740 420 397796 476
rect 396620 364 397796 420
rect 397852 392 398104 476
rect 397880 -960 398104 392
rect 399784 392 400036 480
rect 401660 7924 401716 7934
rect 401660 480 401716 7868
rect 401660 392 401912 480
rect 399784 -960 400008 392
rect 401688 -960 401912 392
rect 403228 420 403284 27692
rect 404908 4788 404964 60060
rect 405468 58828 405524 60060
rect 405020 58772 405524 58828
rect 405020 19348 405076 58772
rect 405020 19282 405076 19292
rect 406588 44548 406644 44558
rect 404908 4722 404964 4732
rect 405468 11172 405524 11182
rect 403452 480 403620 532
rect 405468 480 405524 11116
rect 403452 476 403816 480
rect 403452 420 403508 476
rect 403228 364 403508 420
rect 403564 392 403816 476
rect 405468 392 405720 480
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 406588 420 406644 44492
rect 406700 27860 406756 60060
rect 407372 55524 407428 55534
rect 407372 44548 407428 55468
rect 407372 44482 407428 44492
rect 406700 27794 406756 27804
rect 408268 4676 408324 60060
rect 409948 59106 410004 59118
rect 409948 59054 409950 59106
rect 410002 59054 410004 59106
rect 408268 4610 408324 4620
rect 408380 31108 408436 31118
rect 407260 480 407428 532
rect 407260 476 407624 480
rect 407260 420 407316 476
rect 406588 364 407316 420
rect 407372 392 407624 476
rect 407400 -960 407624 392
rect 408380 420 408436 31052
rect 409948 5908 410004 59054
rect 410060 54852 410116 60060
rect 410732 59106 410788 60060
rect 410732 59054 410734 59106
rect 410786 59054 410788 59106
rect 410732 59042 410788 59054
rect 410060 54786 410116 54796
rect 409948 5842 410004 5852
rect 410060 14308 410116 14318
rect 409164 480 409332 532
rect 409164 476 409528 480
rect 409164 420 409220 476
rect 408380 364 409220 420
rect 409276 392 409528 476
rect 409304 -960 409528 392
rect 410060 420 410116 14252
rect 411628 4564 411684 60060
rect 412412 56756 412468 56766
rect 412412 7700 412468 56700
rect 413308 15988 413364 60060
rect 413308 15922 413364 15932
rect 414988 59442 415044 59454
rect 414988 59390 414990 59442
rect 415042 59390 415044 59442
rect 414988 12740 415044 59390
rect 415100 41300 415156 60088
rect 415660 60060 416360 60116
rect 416668 60060 417592 60116
rect 418348 60060 418824 60116
rect 415660 59442 415716 60060
rect 415660 59390 415662 59442
rect 415714 59390 415716 59442
rect 415660 59378 415716 59390
rect 416668 54740 416724 60060
rect 416668 54674 416724 54684
rect 415100 41234 415156 41244
rect 418348 26068 418404 60060
rect 418348 26002 418404 26012
rect 418460 32900 418516 32910
rect 414988 12674 415044 12684
rect 415772 12628 415828 12638
rect 414988 9380 415044 9390
rect 412412 7634 412468 7644
rect 413084 7812 413140 7822
rect 411628 4498 411684 4508
rect 411068 480 411236 532
rect 413084 480 413140 7756
rect 414988 480 415044 9324
rect 415772 5012 415828 12572
rect 415772 4946 415828 4956
rect 416892 5012 416948 5022
rect 416892 480 416948 4956
rect 411068 476 411432 480
rect 411068 420 411124 476
rect 410060 364 411124 420
rect 411180 392 411432 476
rect 413084 392 413336 480
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418460 420 418516 32844
rect 420028 4452 420084 60088
rect 420140 60060 421288 60116
rect 421820 60060 422520 60116
rect 423388 60060 423752 60116
rect 424060 60060 424984 60116
rect 425068 60060 426216 60116
rect 426748 60060 427448 60116
rect 428428 60060 428680 60116
rect 429100 60060 429912 60116
rect 430108 60060 431144 60116
rect 431788 60060 432376 60116
rect 420140 54628 420196 60060
rect 420140 54562 420196 54572
rect 421708 38052 421764 38062
rect 420028 4386 420084 4396
rect 420700 6244 420756 6254
rect 418684 480 418852 532
rect 420700 480 420756 6188
rect 418684 476 419048 480
rect 418684 420 418740 476
rect 418460 364 418740 420
rect 418796 392 419048 476
rect 420700 392 420952 480
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 421708 420 421764 37996
rect 421820 36148 421876 60060
rect 421820 36082 421876 36092
rect 423388 4340 423444 60060
rect 424060 58828 424116 60060
rect 423500 58772 424116 58828
rect 423500 52948 423556 58772
rect 423500 52882 423556 52892
rect 425068 27748 425124 60060
rect 426748 56868 426804 60060
rect 426748 56802 426804 56812
rect 425068 27682 425124 27692
rect 427532 56308 427588 56318
rect 425068 22820 425124 22830
rect 423388 4274 423444 4284
rect 423500 17892 423556 17902
rect 422492 480 422660 532
rect 422492 476 422856 480
rect 422492 420 422548 476
rect 421708 364 422548 420
rect 422604 392 422856 476
rect 422632 -960 422856 392
rect 423500 420 423556 17836
rect 424396 480 424564 532
rect 424396 476 424760 480
rect 424396 420 424452 476
rect 423500 364 424452 420
rect 424508 392 424760 476
rect 424536 -960 424760 392
rect 425068 420 425124 22764
rect 427532 6804 427588 56252
rect 428428 56308 428484 60060
rect 429100 58828 429156 60060
rect 428428 56242 428484 56252
rect 428540 58772 429156 58828
rect 427532 6738 427588 6748
rect 428428 39508 428484 39518
rect 426300 480 426468 532
rect 428428 480 428484 39452
rect 428540 31108 428596 58772
rect 428540 31042 428596 31052
rect 430108 12628 430164 60060
rect 431788 56756 431844 60060
rect 431788 56690 431844 56700
rect 433468 59444 433524 59454
rect 432572 56532 432628 56542
rect 432572 17892 432628 56476
rect 432572 17826 432628 17836
rect 430108 12562 430164 12572
rect 432124 11060 432180 11070
rect 430220 6804 430276 6814
rect 430220 480 430276 6748
rect 432124 480 432180 11004
rect 433468 4228 433524 59388
rect 433580 14308 433636 60088
rect 434140 60060 434840 60116
rect 434140 59444 434196 60060
rect 434140 59378 434196 59388
rect 436828 21924 436884 438508
rect 440188 41188 440244 442092
rect 441868 438676 441924 438686
rect 440188 41122 440244 41132
rect 440300 46452 440356 46462
rect 436828 21858 436884 21868
rect 433580 14242 433636 14252
rect 436828 21140 436884 21150
rect 433468 4162 433524 4172
rect 433580 12852 433636 12862
rect 426300 476 426664 480
rect 426300 420 426356 476
rect 425068 364 426356 420
rect 426412 392 426664 476
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430220 392 430472 480
rect 432124 392 432376 480
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 433580 420 433636 12796
rect 435932 2660 435988 2670
rect 433916 480 434084 532
rect 435932 480 435988 2604
rect 433916 476 434280 480
rect 433916 420 433972 476
rect 433580 364 433972 420
rect 434028 392 434280 476
rect 435932 392 436184 480
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 436828 420 436884 21084
rect 439740 6132 439796 6142
rect 437724 480 437892 532
rect 439740 480 439796 6076
rect 437724 476 438088 480
rect 437724 420 437780 476
rect 436828 364 437780 420
rect 437836 392 438088 476
rect 439740 392 439992 480
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 440300 420 440356 46396
rect 441868 8484 441924 438620
rect 442652 430164 442708 443996
rect 442652 430098 442708 430108
rect 444332 231924 444388 458892
rect 444332 231858 444388 231868
rect 446012 440580 446068 440590
rect 446012 205044 446068 440524
rect 447692 270564 447748 462140
rect 454412 457828 454468 590492
rect 474348 590548 474404 595560
rect 474348 590482 474404 590492
rect 495628 461300 495684 595644
rect 496300 595476 496356 595644
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 561148 595644 562548 595700
rect 562632 595672 562856 597000
rect 496412 595476 496468 595560
rect 496300 595420 496468 595476
rect 518476 593236 518532 595560
rect 518476 593170 518532 593180
rect 540540 593124 540596 595560
rect 540540 593058 540596 593068
rect 495628 461234 495684 461244
rect 454412 457762 454468 457772
rect 486332 455588 486388 455598
rect 484652 455476 484708 455486
rect 481292 455364 481348 455374
rect 477932 453796 477988 453806
rect 476252 452116 476308 452126
rect 466172 450772 466228 450782
rect 464492 450548 464548 450558
rect 459452 450324 459508 450334
rect 456092 445508 456148 445518
rect 451052 443828 451108 443838
rect 449372 442036 449428 442046
rect 449372 416724 449428 441980
rect 449372 416658 449428 416668
rect 451052 362964 451108 443772
rect 451052 362898 451108 362908
rect 454412 441924 454468 441934
rect 447692 270498 447748 270508
rect 446012 204978 446068 204988
rect 454412 178164 454468 441868
rect 454412 178098 454468 178108
rect 456092 112644 456148 445452
rect 459452 218484 459508 450268
rect 464492 310884 464548 450492
rect 466172 349524 466228 450716
rect 467852 445620 467908 445630
rect 467852 389844 467908 445564
rect 467852 389778 467908 389788
rect 466172 349458 466228 349468
rect 464492 310818 464548 310828
rect 459452 218418 459508 218428
rect 456092 112578 456148 112588
rect 476252 99204 476308 452060
rect 477932 137844 477988 453740
rect 479612 447300 479668 447310
rect 479612 257124 479668 447244
rect 481292 297444 481348 455308
rect 484652 336084 484708 455420
rect 486332 376404 486388 455532
rect 487788 455364 487844 455374
rect 487788 454468 487844 455308
rect 487788 454402 487844 454412
rect 486332 376338 486388 376348
rect 496412 447076 496468 447086
rect 484652 336018 484708 336028
rect 481292 297378 481348 297388
rect 479612 257058 479668 257068
rect 477932 137778 477988 137788
rect 476252 99138 476308 99148
rect 496412 58884 496468 447020
rect 561148 442708 561204 595644
rect 562492 595476 562548 595644
rect 562604 595560 562856 595672
rect 584696 595672 584920 597000
rect 584696 595560 584948 595672
rect 562604 595476 562660 595560
rect 562492 595420 562660 595476
rect 584892 590548 584948 595560
rect 584892 590482 584948 590492
rect 593292 590548 593348 590558
rect 593068 562212 593124 562222
rect 593068 464548 593124 562156
rect 593180 522564 593236 522574
rect 593180 466228 593236 522508
rect 593292 467908 593348 590492
rect 593292 467842 593348 467852
rect 593740 473844 593796 473854
rect 593180 466162 593236 466172
rect 593404 467124 593460 467134
rect 593068 464482 593124 464492
rect 593180 465444 593236 465454
rect 590492 448644 590548 448654
rect 588812 446964 588868 446984
rect 588812 443492 588868 446908
rect 588812 443426 588868 443436
rect 561148 442642 561204 442652
rect 590492 192388 590548 448588
rect 593068 440244 593124 440254
rect 593068 403844 593124 440188
rect 593068 403778 593124 403788
rect 590492 192322 590548 192332
rect 496412 58818 496468 58828
rect 458668 58100 458724 58110
rect 446012 56868 446068 56878
rect 444332 56644 444388 56654
rect 441868 8418 441924 8428
rect 443548 17780 443604 17790
rect 441532 480 441700 532
rect 443548 480 443604 17724
rect 444332 9380 444388 56588
rect 446012 39508 446068 56812
rect 454412 56756 454468 56766
rect 448588 54964 448644 54974
rect 446012 39442 446068 39452
rect 446908 44772 446964 44782
rect 445228 34580 445284 34590
rect 445228 11788 445284 34524
rect 445228 11732 445508 11788
rect 444332 9314 444388 9324
rect 445452 480 445508 11732
rect 441532 476 441896 480
rect 441532 420 441588 476
rect 440300 364 441588 420
rect 441644 392 441896 476
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 446908 420 446964 44716
rect 447244 480 447412 532
rect 447244 476 447608 480
rect 447244 420 447300 476
rect 446908 364 447300 420
rect 447356 392 447608 476
rect 447384 -960 447608 392
rect 448588 420 448644 54908
rect 450268 53172 450324 53182
rect 449148 480 449316 532
rect 449148 476 449512 480
rect 449148 420 449204 476
rect 448588 364 449204 420
rect 449260 392 449512 476
rect 449288 -960 449512 392
rect 450268 420 450324 53116
rect 454412 32900 454468 56700
rect 454412 32834 454468 32844
rect 453628 29540 453684 29550
rect 451948 16100 452004 16110
rect 451052 480 451220 532
rect 451052 476 451416 480
rect 451052 420 451108 476
rect 450268 364 451108 420
rect 451164 392 451416 476
rect 451192 -960 451416 392
rect 451948 420 452004 16044
rect 452956 480 453124 532
rect 452956 476 453320 480
rect 452956 420 453012 476
rect 451948 364 453012 420
rect 453068 392 453320 476
rect 453096 -960 453320 392
rect 453628 420 453684 29484
rect 456092 19460 456148 19470
rect 456092 5012 456148 19404
rect 458668 11788 458724 58044
rect 493948 57988 494004 57998
rect 484652 56420 484708 56430
rect 465388 51492 465444 51502
rect 462028 48132 462084 48142
rect 460348 36260 460404 36270
rect 458668 11732 458836 11788
rect 456092 4946 456148 4956
rect 456988 5012 457044 5022
rect 454860 480 455028 532
rect 456988 480 457044 4956
rect 458780 480 458836 11732
rect 454860 476 455224 480
rect 454860 420 454916 476
rect 453628 364 454916 420
rect 454972 392 455224 476
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 458808 -960 459032 392
rect 460348 420 460404 36204
rect 460572 480 460740 532
rect 460572 476 460936 480
rect 460572 420 460628 476
rect 460348 364 460628 420
rect 460684 392 460936 476
rect 460712 -960 460936 392
rect 462028 420 462084 48076
rect 463708 41412 463764 41422
rect 462476 480 462644 532
rect 462476 476 462840 480
rect 462476 420 462532 476
rect 462028 364 462532 420
rect 462588 392 462840 476
rect 462616 -960 462840 392
rect 463708 420 463764 41356
rect 464380 480 464548 532
rect 464380 476 464744 480
rect 464380 420 464436 476
rect 463708 364 464436 420
rect 464492 392 464744 476
rect 464520 -960 464744 392
rect 465388 420 465444 51436
rect 472108 51380 472164 51390
rect 467068 39620 467124 39630
rect 466284 480 466452 532
rect 466284 476 466648 480
rect 466284 420 466340 476
rect 465388 364 466340 420
rect 466396 392 466648 476
rect 466424 -960 466648 392
rect 467068 420 467124 39564
rect 468748 21028 468804 21038
rect 468188 480 468356 532
rect 468188 476 468552 480
rect 468188 420 468244 476
rect 467068 364 468244 420
rect 468300 392 468552 476
rect 468328 -960 468552 392
rect 468748 420 468804 20972
rect 470092 480 470260 532
rect 472108 480 472164 51324
rect 480508 46340 480564 46350
rect 477148 42980 477204 42990
rect 475468 17892 475524 17902
rect 474012 6020 474068 6030
rect 474012 480 474068 5964
rect 470092 476 470456 480
rect 470092 420 470148 476
rect 468748 364 470148 420
rect 470204 392 470456 476
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475468 420 475524 17836
rect 475804 480 475972 532
rect 475804 476 476168 480
rect 475804 420 475860 476
rect 475468 364 475860 420
rect 475916 392 476168 476
rect 475944 -960 476168 392
rect 477148 420 477204 42924
rect 478828 26180 478884 26190
rect 477708 480 477876 532
rect 477708 476 478072 480
rect 477708 420 477764 476
rect 477148 364 477764 420
rect 477820 392 478072 476
rect 477848 -960 478072 392
rect 478828 420 478884 26124
rect 479612 480 479780 532
rect 479612 476 479976 480
rect 479612 420 479668 476
rect 478828 364 479668 420
rect 479724 392 479976 476
rect 479752 -960 479976 392
rect 480508 420 480564 46284
rect 482188 29428 482244 29438
rect 481516 480 481684 532
rect 481516 476 481880 480
rect 481516 420 481572 476
rect 480508 364 481572 420
rect 481628 392 481880 476
rect 481656 -960 481880 392
rect 482188 420 482244 29372
rect 484652 6020 484708 56364
rect 487228 53060 487284 53070
rect 484652 5954 484708 5964
rect 485548 31220 485604 31230
rect 483420 480 483588 532
rect 485548 480 485604 31164
rect 487228 11788 487284 53004
rect 490588 34468 490644 34478
rect 487228 11732 487396 11788
rect 487340 480 487396 11732
rect 489244 7588 489300 7598
rect 489244 480 489300 7532
rect 483420 476 483784 480
rect 483420 420 483476 476
rect 482188 364 483476 420
rect 483532 392 483784 476
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 490588 420 490644 34412
rect 493052 2548 493108 2558
rect 491036 480 491204 532
rect 493052 480 493108 2492
rect 491036 476 491400 480
rect 491036 420 491092 476
rect 490588 364 491092 420
rect 491148 392 491400 476
rect 493052 392 493304 480
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 493948 420 494004 57932
rect 570332 56308 570388 56318
rect 544348 54852 544404 54862
rect 522508 51268 522564 51278
rect 505708 49700 505764 49710
rect 502348 48020 502404 48030
rect 500668 46228 500724 46238
rect 497308 22708 497364 22718
rect 496860 9268 496916 9278
rect 494844 480 495012 532
rect 496860 480 496916 9212
rect 494844 476 495208 480
rect 494844 420 494900 476
rect 493948 364 494900 420
rect 494956 392 495208 476
rect 496860 392 497112 480
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 497308 420 497364 22652
rect 498652 480 498820 532
rect 500668 480 500724 46172
rect 502348 11788 502404 47964
rect 504028 24500 504084 24510
rect 502348 11732 502628 11788
rect 502572 480 502628 11732
rect 498652 476 499016 480
rect 498652 420 498708 476
rect 497308 364 498708 420
rect 498764 392 499016 476
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504028 420 504084 24444
rect 504364 480 504532 532
rect 504364 476 504728 480
rect 504364 420 504420 476
rect 504028 364 504420 420
rect 504476 392 504728 476
rect 504504 -960 504728 392
rect 505708 420 505764 49644
rect 514108 47908 514164 47918
rect 512428 37940 512484 37950
rect 509068 24388 509124 24398
rect 508284 6020 508340 6030
rect 506268 480 506436 532
rect 508284 480 508340 5964
rect 506268 476 506632 480
rect 506268 420 506324 476
rect 505708 364 506324 420
rect 506380 392 506632 476
rect 508284 392 508536 480
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 509068 420 509124 24332
rect 512428 5012 512484 37884
rect 512316 4956 512484 5012
rect 510076 480 510244 532
rect 512316 480 512372 4956
rect 514108 480 514164 47852
rect 515788 44660 515844 44670
rect 515788 11788 515844 44604
rect 520828 32788 520884 32798
rect 515788 11732 515956 11788
rect 515900 480 515956 11732
rect 517804 10948 517860 10958
rect 517804 480 517860 10892
rect 519708 7700 519764 7710
rect 519708 480 519764 7644
rect 510076 476 510440 480
rect 510076 420 510132 476
rect 509068 364 510132 420
rect 510188 392 510440 476
rect 510216 -960 510440 392
rect 512120 392 512372 480
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 520828 420 520884 32732
rect 521500 480 521668 532
rect 521500 476 521864 480
rect 521500 420 521556 476
rect 520828 364 521556 420
rect 521612 392 521864 476
rect 521640 -960 521864 392
rect 522508 420 522564 51212
rect 534268 49588 534324 49598
rect 530908 44548 530964 44558
rect 523292 17668 523348 17678
rect 523292 5012 523348 17612
rect 529228 14420 529284 14430
rect 527324 9380 527380 9390
rect 523292 4946 523348 4956
rect 525420 5012 525476 5022
rect 523404 480 523572 532
rect 525420 480 525476 4956
rect 527324 480 527380 9324
rect 529228 480 529284 14364
rect 530908 11788 530964 44492
rect 532588 37828 532644 37838
rect 530908 11732 531188 11788
rect 531132 480 531188 11732
rect 523404 476 523768 480
rect 523404 420 523460 476
rect 522508 364 523460 420
rect 523516 392 523768 476
rect 525420 392 525672 480
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 532588 420 532644 37772
rect 532924 480 533092 532
rect 532924 476 533288 480
rect 532924 420 532980 476
rect 532588 364 532980 420
rect 533036 392 533288 476
rect 533064 -960 533288 392
rect 534268 420 534324 49532
rect 539308 27860 539364 27870
rect 537628 19348 537684 19358
rect 536844 4788 536900 4798
rect 534828 480 534996 532
rect 536844 480 536900 4732
rect 534828 476 535192 480
rect 534828 420 534884 476
rect 534268 364 534884 420
rect 534940 392 535192 476
rect 536844 392 537096 480
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 537628 420 537684 19292
rect 538636 480 538804 532
rect 538636 476 539000 480
rect 538636 420 538692 476
rect 537628 364 538692 420
rect 538748 392 539000 476
rect 538776 -960 539000 392
rect 539308 420 539364 27804
rect 544348 11788 544404 54796
rect 554428 54740 554484 54750
rect 551068 41300 551124 41310
rect 549388 15988 549444 15998
rect 544348 11732 544516 11788
rect 542668 4676 542724 4686
rect 540540 480 540708 532
rect 542668 480 542724 4620
rect 544460 480 544516 11732
rect 546364 5908 546420 5918
rect 546364 480 546420 5852
rect 548268 4564 548324 4574
rect 548268 480 548324 4508
rect 540540 476 540904 480
rect 540540 420 540596 476
rect 539308 364 540596 420
rect 540652 392 540904 476
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 549388 420 549444 15932
rect 550060 480 550228 532
rect 550060 476 550424 480
rect 550060 420 550116 476
rect 549388 364 550116 420
rect 550172 392 550424 476
rect 550200 -960 550424 392
rect 551068 420 551124 41244
rect 552748 12740 552804 12750
rect 551964 480 552132 532
rect 551964 476 552328 480
rect 551964 420 552020 476
rect 551068 364 552020 420
rect 552076 392 552328 476
rect 552104 -960 552328 392
rect 552748 420 552804 12684
rect 553868 480 554036 532
rect 553868 476 554232 480
rect 553868 420 553924 476
rect 552748 364 553924 420
rect 553980 392 554232 476
rect 554008 -960 554232 392
rect 554428 420 554484 54684
rect 560252 54628 560308 54638
rect 557788 26068 557844 26078
rect 555772 480 555940 532
rect 557788 480 557844 26012
rect 560252 5012 560308 54572
rect 566188 52948 566244 52958
rect 562828 36148 562884 36158
rect 560252 4946 560308 4956
rect 561596 5012 561652 5022
rect 559692 4452 559748 4462
rect 559692 480 559748 4396
rect 561596 480 561652 4956
rect 555772 476 556136 480
rect 555772 420 555828 476
rect 554428 364 555828 420
rect 555884 392 556136 476
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 562828 420 562884 36092
rect 565404 4340 565460 4350
rect 563388 480 563556 532
rect 565404 480 565460 4284
rect 563388 476 563752 480
rect 563388 420 563444 476
rect 562828 364 563444 420
rect 563500 392 563752 476
rect 565404 392 565656 480
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 566188 420 566244 52892
rect 567868 27748 567924 27758
rect 567196 480 567364 532
rect 567196 476 567560 480
rect 567196 420 567252 476
rect 566188 364 567252 420
rect 567308 392 567560 476
rect 567336 -960 567560 392
rect 567868 420 567924 27692
rect 570332 10164 570388 56252
rect 590492 42868 590548 42878
rect 570332 10098 570388 10108
rect 571228 39508 571284 39518
rect 569100 480 569268 532
rect 571228 480 571284 39452
rect 579628 32900 579684 32910
rect 574588 31108 574644 31118
rect 573020 10164 573076 10174
rect 573020 480 573076 10108
rect 569100 476 569464 480
rect 569100 420 569156 476
rect 567868 364 569156 420
rect 569212 392 569464 476
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 573048 -960 573272 392
rect 574588 420 574644 31052
rect 576268 12628 576324 12638
rect 574812 480 574980 532
rect 574812 476 575176 480
rect 574812 420 574868 476
rect 574588 364 574868 420
rect 574924 392 575176 476
rect 574952 -960 575176 392
rect 576268 420 576324 12572
rect 576716 480 576884 532
rect 576716 476 577080 480
rect 576716 420 576772 476
rect 576268 364 576772 420
rect 576828 392 577080 476
rect 576856 -960 577080 392
rect 578760 -960 578984 480
rect 579628 420 579684 32844
rect 590492 20580 590548 42812
rect 593180 33796 593236 465388
rect 593292 445284 593348 445294
rect 593292 47012 593348 445228
rect 593404 73444 593460 467068
rect 593628 458724 593684 458734
rect 593516 457044 593572 457054
rect 593516 86660 593572 456988
rect 593628 126308 593684 458668
rect 593740 152740 593796 473788
rect 594076 470484 594132 470504
rect 593852 462084 593908 462094
rect 593852 165956 593908 462028
rect 593964 452004 594020 452014
rect 593964 245252 594020 451948
rect 594076 284900 594132 470428
rect 594188 460404 594244 460414
rect 594188 324548 594244 460348
rect 594188 324482 594244 324492
rect 594300 443604 594356 443614
rect 594076 284834 594132 284844
rect 593964 245186 594020 245196
rect 593852 165890 593908 165900
rect 593740 152674 593796 152684
rect 593628 126242 593684 126252
rect 593516 86594 593572 86604
rect 593404 73378 593460 73388
rect 593292 46946 593348 46956
rect 593180 33730 593236 33740
rect 590492 20514 590548 20524
rect 581308 14308 581364 14318
rect 580524 480 580692 532
rect 580524 476 580888 480
rect 580524 420 580580 476
rect 579628 364 580580 420
rect 580636 392 580888 476
rect 580664 -960 580888 392
rect 581308 420 581364 14252
rect 594300 7364 594356 443548
rect 594300 7298 594356 7308
rect 584444 4228 584500 4238
rect 582428 480 582596 532
rect 584444 480 584500 4172
rect 582428 476 582792 480
rect 582428 420 582484 476
rect 581308 364 582484 420
rect 582540 392 582792 476
rect 584444 392 584696 480
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 5852 530684 5908 530740
rect 4172 516572 4228 516628
rect 2492 468860 2548 468916
rect 5852 462812 5908 462868
rect 9212 463708 9268 463764
rect 4172 442764 4228 442820
rect 5852 447132 5908 447188
rect 5852 291004 5908 291060
rect 55356 593292 55412 593348
rect 33292 590492 33348 590548
rect 12572 557788 12628 557844
rect 14252 473788 14308 473844
rect 14252 461132 14308 461188
rect 17612 472108 17668 472164
rect 12572 459452 12628 459508
rect 15932 457100 15988 457156
rect 14252 455644 14308 455700
rect 10108 442876 10164 442932
rect 12572 443660 12628 443716
rect 10892 438508 10948 438564
rect 14252 431788 14308 431844
rect 12572 332668 12628 332724
rect 15932 304108 15988 304164
rect 10892 220444 10948 220500
rect 9212 121660 9268 121716
rect 2492 107436 2548 107492
rect 22652 470540 22708 470596
rect 19292 465500 19348 465556
rect 19292 317548 19348 317604
rect 22652 191548 22708 191604
rect 27692 467180 27748 467236
rect 68908 465388 68964 465444
rect 36092 463820 36148 463876
rect 31052 452284 31108 452340
rect 29372 448812 29428 448868
rect 31052 361228 31108 361284
rect 32732 448700 32788 448756
rect 29372 176428 29428 176484
rect 27692 149548 27748 149604
rect 32732 134428 32788 134484
rect 34412 440300 34468 440356
rect 17612 92428 17668 92484
rect 28588 56252 28644 56308
rect 4956 41132 5012 41188
rect 4956 36876 5012 36932
rect 19292 36204 19348 36260
rect 15148 36092 15204 36148
rect 10108 22652 10164 22708
rect 13356 5852 13412 5908
rect 17276 4956 17332 5012
rect 27692 12684 27748 12740
rect 19292 4956 19348 5012
rect 22988 10892 23044 10948
rect 21084 4284 21140 4340
rect 19180 4172 19236 4228
rect 24892 4956 24948 5012
rect 27692 4956 27748 5012
rect 26796 4844 26852 4900
rect 31948 52892 32004 52948
rect 30268 20972 30324 21028
rect 52892 453852 52948 453908
rect 44492 453628 44548 453684
rect 41132 452172 41188 452228
rect 37772 450380 37828 450436
rect 37772 275548 37828 275604
rect 36092 262108 36148 262164
rect 41132 233548 41188 233604
rect 44604 449036 44660 449092
rect 51212 448924 51268 448980
rect 44604 403228 44660 403284
rect 46172 447356 46228 447412
rect 47852 445676 47908 445732
rect 47852 388108 47908 388164
rect 49532 440412 49588 440468
rect 46172 346108 46228 346164
rect 54572 450604 54628 450660
rect 56252 443884 56308 443940
rect 66444 443548 66500 443604
rect 60396 441868 60452 441924
rect 59612 440636 59668 440692
rect 59612 416668 59668 416724
rect 56252 374668 56308 374724
rect 54572 246988 54628 247044
rect 52892 204988 52948 205044
rect 51212 162988 51268 163044
rect 49532 78988 49588 79044
rect 44492 63868 44548 63924
rect 56252 56364 56308 56420
rect 53788 54796 53844 54852
rect 36092 54684 36148 54740
rect 34412 50428 34468 50484
rect 34524 53004 34580 53060
rect 34524 4844 34580 4900
rect 34412 4508 34468 4564
rect 36988 54572 37044 54628
rect 36092 4508 36148 4564
rect 36316 7532 36372 7588
rect 40348 51212 40404 51268
rect 40124 4956 40180 5012
rect 44492 27692 44548 27748
rect 48748 26012 48804 26068
rect 47068 19292 47124 19348
rect 45388 17612 45444 17668
rect 44492 4956 44548 5012
rect 43932 4396 43988 4452
rect 52108 25116 52164 25172
rect 51548 4508 51604 4564
rect 56252 25116 56308 25172
rect 58828 44492 58884 44548
rect 76188 445228 76244 445284
rect 72940 441868 72996 441924
rect 99484 591276 99540 591332
rect 104972 591276 105028 591332
rect 97468 473788 97524 473844
rect 77308 442988 77364 443044
rect 78988 467068 79044 467124
rect 94108 458668 94164 458724
rect 85708 456988 85764 457044
rect 82348 447020 82404 447076
rect 92428 452060 92484 452116
rect 89180 445452 89236 445508
rect 104188 462028 104244 462084
rect 100828 453740 100884 453796
rect 120988 474572 121044 474628
rect 134428 470428 134484 470484
rect 104972 461356 105028 461412
rect 127708 462140 127764 462196
rect 117628 458892 117684 458948
rect 108668 442652 108724 442708
rect 111916 441868 111972 441924
rect 115164 440524 115220 440580
rect 124348 451948 124404 452004
rect 120988 450268 121044 450324
rect 131068 447244 131124 447300
rect 142828 457996 142884 458052
rect 142940 460348 142996 460404
rect 141148 455308 141204 455364
rect 137788 450492 137844 450548
rect 159628 455532 159684 455588
rect 149548 455420 149604 455476
rect 146188 450716 146244 450772
rect 157388 445564 157444 445620
rect 154140 443772 154196 443828
rect 187740 590604 187796 590660
rect 188972 590604 189028 590660
rect 185612 482188 185668 482244
rect 176428 468748 176484 468804
rect 170492 448588 170548 448644
rect 164668 443100 164724 443156
rect 167132 443996 167188 444052
rect 163884 440188 163940 440244
rect 170492 442652 170548 442708
rect 173068 446908 173124 446964
rect 170380 441980 170436 442036
rect 179788 454412 179844 454468
rect 183372 444108 183428 444164
rect 207452 588028 207508 588084
rect 194908 547708 194964 547764
rect 194012 509068 194068 509124
rect 188972 472892 189028 472948
rect 189868 495628 189924 495684
rect 185612 444108 185668 444164
rect 186620 444332 186676 444388
rect 191548 466172 191604 466228
rect 198268 534268 198324 534324
rect 201628 464492 201684 464548
rect 194012 444332 194068 444388
rect 206108 444108 206164 444164
rect 224252 593180 224308 593236
rect 208572 575372 208628 575428
rect 215068 593068 215124 593124
rect 208348 574588 208404 574644
rect 212492 502348 212548 502404
rect 212492 476252 212548 476308
rect 211708 467852 211764 467908
rect 207452 444108 207508 444164
rect 222348 443212 222404 443268
rect 219100 442652 219156 442708
rect 230188 464604 230244 464660
rect 231868 593404 231924 593460
rect 228508 461244 228564 461300
rect 224252 443212 224308 443268
rect 225148 457772 225204 457828
rect 242732 590604 242788 590660
rect 238588 469532 238644 469588
rect 235228 457884 235284 457940
rect 241836 444108 241892 444164
rect 250348 503132 250404 503188
rect 246988 462924 247044 462980
rect 243628 459564 243684 459620
rect 246092 458780 246148 458836
rect 246092 454524 246148 454580
rect 274652 590492 274708 590548
rect 263788 575372 263844 575428
rect 253708 471212 253764 471268
rect 260428 471212 260484 471268
rect 257068 463036 257124 463092
rect 253708 459676 253764 459732
rect 242732 444108 242788 444164
rect 270508 472892 270564 472948
rect 267148 464604 267204 464660
rect 273868 457996 273924 458052
rect 288988 593292 289044 593348
rect 275548 459676 275604 459732
rect 280588 474572 280644 474628
rect 274652 457996 274708 458052
rect 277564 443100 277620 443156
rect 287308 461356 287364 461412
rect 284060 442988 284116 443044
rect 303212 590492 303268 590548
rect 297388 463036 297444 463092
rect 299068 586348 299124 586404
rect 295708 457996 295764 458052
rect 303212 462924 303268 462980
rect 305788 572908 305844 572964
rect 302428 459452 302484 459508
rect 308252 544348 308308 544404
rect 293804 442876 293860 442932
rect 319228 503132 319284 503188
rect 325052 487228 325108 487284
rect 319228 476252 319284 476308
rect 315868 462812 315924 462868
rect 308252 443100 308308 443156
rect 310044 443100 310100 443156
rect 313292 442764 313348 442820
rect 322588 461132 322644 461188
rect 386092 590604 386148 590660
rect 364028 590492 364084 590548
rect 393148 470540 393204 470596
rect 341068 459564 341124 459620
rect 364588 465500 364644 465556
rect 361228 457100 361284 457156
rect 332668 455644 332724 455700
rect 329308 454524 329364 454580
rect 325052 448476 325108 448532
rect 325948 448476 326004 448532
rect 354508 452284 354564 452340
rect 344428 449036 344484 449092
rect 351148 447356 351204 447412
rect 342524 445676 342580 445732
rect 336028 445340 336084 445396
rect 339276 440636 339332 440692
rect 349020 443884 349076 443940
rect 358764 443660 358820 443716
rect 371308 463820 371364 463876
rect 367948 447132 368004 447188
rect 386428 453852 386484 453908
rect 384748 452172 384804 452228
rect 378028 450604 378084 450660
rect 374668 450380 374724 450436
rect 389788 448812 389844 448868
rect 403228 467180 403284 467236
rect 396508 448924 396564 448980
rect 399868 448700 399924 448756
rect 406588 463708 406644 463764
rect 427532 590828 427588 590884
rect 408268 457884 408324 457940
rect 409948 472108 410004 472164
rect 451612 593404 451668 593460
rect 430220 590828 430276 590884
rect 427532 469532 427588 469588
rect 454412 590492 454468 590548
rect 413308 468860 413364 468916
rect 447692 462140 447748 462196
rect 444332 458892 444388 458948
rect 423388 453628 423444 453684
rect 417228 440412 417284 440468
rect 420476 440300 420532 440356
rect 442652 443996 442708 444052
rect 426972 442092 427028 442148
rect 440188 442092 440244 442148
rect 381500 439292 381556 439348
rect 430220 439292 430276 439348
rect 433468 439292 433524 439348
rect 436828 438508 436884 438564
rect 60396 42812 60452 42868
rect 62972 56588 63028 56644
rect 57260 4620 57316 4676
rect 63868 22652 63924 22708
rect 62972 10892 63028 10948
rect 63868 15932 63924 15988
rect 61068 5964 61124 6020
rect 62972 4732 63028 4788
rect 67228 36092 67284 36148
rect 68012 56476 68068 56532
rect 68012 5964 68068 6020
rect 65548 5852 65604 5908
rect 66780 5852 66836 5908
rect 68684 4844 68740 4900
rect 69020 36204 69076 36260
rect 68908 4172 68964 4228
rect 69020 14252 69076 14308
rect 72268 56588 72324 56644
rect 75628 56252 75684 56308
rect 73948 53004 74004 53060
rect 76412 55468 76468 55524
rect 77308 55468 77364 55524
rect 76412 20972 76468 21028
rect 77308 53116 77364 53172
rect 72716 12684 72772 12740
rect 75628 16044 75684 16100
rect 70588 4284 70644 4340
rect 72492 12572 72548 12628
rect 74396 4172 74452 4228
rect 78988 54684 79044 54740
rect 77420 52892 77476 52948
rect 82460 54572 82516 54628
rect 83132 56588 83188 56644
rect 82348 27692 82404 27748
rect 82348 20972 82404 21028
rect 80668 7532 80724 7588
rect 82012 7756 82068 7812
rect 80108 4284 80164 4340
rect 84028 51212 84084 51268
rect 84812 55468 84868 55524
rect 84812 17612 84868 17668
rect 83132 5852 83188 5908
rect 82908 4956 82964 5012
rect 82908 4508 82964 4564
rect 87388 55468 87444 55524
rect 90748 59388 90804 59444
rect 90748 56364 90804 56420
rect 89180 55468 89236 55524
rect 89180 54796 89236 54852
rect 89068 26012 89124 26068
rect 87500 19292 87556 19348
rect 89628 10892 89684 10948
rect 85708 4508 85764 4564
rect 87724 5852 87780 5908
rect 85820 4396 85876 4452
rect 91644 59388 91700 59444
rect 91532 56700 91588 56756
rect 92428 55468 92484 55524
rect 91532 44492 91588 44548
rect 90972 4956 91028 5012
rect 91532 6076 91588 6132
rect 93436 5964 93492 6020
rect 95788 56700 95844 56756
rect 95900 56476 95956 56532
rect 94892 56252 94948 56308
rect 94892 6076 94948 6132
rect 95340 7532 95396 7588
rect 94108 4620 94164 4676
rect 98700 56700 98756 56756
rect 98700 53116 98756 53172
rect 100828 56588 100884 56644
rect 99148 15932 99204 15988
rect 99932 56476 99988 56532
rect 99932 7756 99988 7812
rect 97468 4732 97524 4788
rect 99036 7644 99092 7700
rect 97244 4508 97300 4564
rect 102508 14252 102564 14308
rect 102732 14252 102788 14308
rect 100940 4844 100996 4900
rect 101052 4620 101108 4676
rect 104188 12572 104244 12628
rect 104412 12572 104468 12628
rect 107548 56700 107604 56756
rect 109228 59388 109284 59444
rect 109228 56476 109284 56532
rect 105980 16044 106036 16100
rect 107548 56364 107604 56420
rect 105868 4172 105924 4228
rect 106764 4172 106820 4228
rect 110124 59388 110180 59444
rect 110012 55468 110068 55524
rect 110908 55468 110964 55524
rect 110012 20972 110068 21028
rect 109452 4284 109508 4340
rect 110572 6076 110628 6132
rect 114268 59388 114324 59444
rect 113372 55468 113428 55524
rect 114268 55468 114324 55524
rect 115052 59388 115108 59444
rect 115948 56252 116004 56308
rect 114492 55468 114548 55524
rect 116060 55468 116116 55524
rect 113372 10892 113428 10948
rect 115948 15932 116004 15988
rect 118412 55468 118468 55524
rect 119308 55468 119364 55524
rect 118412 7532 118468 7588
rect 117628 5964 117684 6020
rect 112588 4396 112644 4452
rect 114380 4396 114436 4452
rect 112476 4284 112532 4340
rect 116172 5852 116228 5908
rect 118188 4732 118244 4788
rect 119532 4508 119588 4564
rect 120092 9212 120148 9268
rect 120988 7644 121044 7700
rect 121996 7532 122052 7588
rect 123452 55468 123508 55524
rect 124348 55468 124404 55524
rect 124460 14252 124516 14308
rect 125132 56252 125188 56308
rect 123452 12572 123508 12628
rect 122668 4620 122724 4676
rect 123900 5852 123956 5908
rect 125132 5852 125188 5908
rect 125804 5852 125860 5908
rect 127708 56364 127764 56420
rect 128492 56364 128548 56420
rect 128492 15932 128548 15988
rect 127820 6076 127876 6132
rect 126028 4172 126084 4228
rect 127596 5964 127652 6020
rect 132748 56364 132804 56420
rect 131852 55468 131908 55524
rect 131852 9212 131908 9268
rect 131068 4396 131124 4452
rect 132636 7644 132692 7700
rect 129388 4284 129444 4340
rect 131516 3836 131572 3892
rect 129612 3388 129668 3444
rect 134428 55468 134484 55524
rect 135212 56476 135268 56532
rect 132860 4732 132916 4788
rect 133420 4956 133476 5012
rect 132636 3388 132692 3444
rect 135436 55468 135492 55524
rect 136108 55468 136164 55524
rect 136220 56364 136276 56420
rect 137788 56252 137844 56308
rect 135436 7532 135492 7588
rect 135212 4956 135268 5012
rect 135324 4172 135380 4228
rect 137788 7532 137844 7588
rect 139468 5964 139524 6020
rect 140252 56588 140308 56644
rect 137900 5852 137956 5908
rect 137788 3836 137844 3892
rect 139132 4956 139188 5012
rect 142828 59388 142884 59444
rect 142828 56476 142884 56532
rect 141148 7644 141204 7700
rect 142716 7980 142772 8036
rect 140252 4956 140308 5012
rect 141036 5852 141092 5908
rect 143388 59388 143444 59444
rect 143276 7532 143332 7588
rect 144508 55580 144564 55636
rect 142716 4172 142772 4228
rect 142940 6748 142996 6804
rect 146188 59388 146244 59444
rect 146188 56588 146244 56644
rect 147084 59388 147140 59444
rect 146300 56364 146356 56420
rect 144732 7980 144788 8036
rect 147868 5852 147924 5908
rect 148652 55468 148708 55524
rect 146748 4956 146804 5012
rect 151340 55580 151396 55636
rect 151228 55468 151284 55524
rect 149548 6748 149604 6804
rect 152460 7532 152516 7588
rect 148652 4956 148708 5012
rect 150556 4284 150612 4340
rect 148652 4172 148708 4228
rect 152908 4172 152964 4228
rect 154364 4956 154420 5012
rect 156380 7532 156436 7588
rect 156268 4956 156324 5012
rect 154588 4284 154644 4340
rect 156156 4844 156212 4900
rect 157948 4844 158004 4900
rect 158172 4956 158228 5012
rect 159628 4956 159684 5012
rect 160076 4956 160132 5012
rect 161420 4956 161476 5012
rect 164780 55468 164836 55524
rect 166348 4956 166404 5012
rect 166460 55468 166516 55524
rect 168028 55468 168084 55524
rect 169372 4956 169428 5012
rect 169708 4956 169764 5012
rect 171612 56364 171668 56420
rect 169932 4844 169988 4900
rect 171388 55468 171444 55524
rect 173068 4396 173124 4452
rect 173180 4956 173236 5012
rect 174860 56252 174916 56308
rect 176428 56364 176484 56420
rect 174748 4508 174804 4564
rect 175084 4844 175140 4900
rect 176652 55468 176708 55524
rect 178892 55468 178948 55524
rect 178892 4844 178948 4900
rect 178108 4172 178164 4228
rect 178892 4396 178948 4452
rect 179900 5852 179956 5908
rect 180572 56252 180628 56308
rect 181468 7532 181524 7588
rect 180572 4956 180628 5012
rect 182700 4956 182756 5012
rect 179788 4284 179844 4340
rect 180796 4508 180852 4564
rect 184828 56252 184884 56308
rect 183260 55468 183316 55524
rect 185612 55468 185668 55524
rect 185612 6188 185668 6244
rect 183148 4956 183204 5012
rect 184604 4844 184660 4900
rect 188188 4844 188244 4900
rect 186508 4508 186564 4564
rect 190652 56252 190708 56308
rect 190652 6300 190708 6356
rect 189868 4620 189924 4676
rect 190316 5852 190372 5908
rect 188524 4396 188580 4452
rect 188412 4284 188468 4340
rect 186508 4172 186564 4228
rect 193228 59388 193284 59444
rect 191548 4284 191604 4340
rect 192220 7532 192276 7588
rect 193900 59388 193956 59444
rect 199948 55580 200004 55636
rect 198380 12684 198436 12740
rect 198268 10892 198324 10948
rect 196588 7756 196644 7812
rect 197932 6300 197988 6356
rect 194908 5964 194964 6020
rect 196028 6188 196084 6244
rect 193452 4732 193508 4788
rect 194124 4956 194180 5012
rect 193228 4172 193284 4228
rect 199948 4508 200004 4564
rect 203308 56476 203364 56532
rect 201740 55468 201796 55524
rect 202412 55580 202468 55636
rect 202412 14252 202468 14308
rect 204092 55468 204148 55524
rect 204092 7532 204148 7588
rect 201628 4508 201684 4564
rect 201740 4844 201796 4900
rect 203644 4396 203700 4452
rect 206780 55468 206836 55524
rect 206668 5852 206724 5908
rect 204988 4396 205044 4452
rect 205548 4620 205604 4676
rect 207452 4284 207508 4340
rect 210028 56364 210084 56420
rect 210812 56476 210868 56532
rect 209132 55468 209188 55524
rect 209132 16156 209188 16212
rect 210812 6076 210868 6132
rect 208348 4284 208404 4340
rect 209356 4732 209412 4788
rect 211260 4172 211316 4228
rect 211820 56476 211876 56532
rect 213388 56252 213444 56308
rect 214172 56364 214228 56420
rect 215068 12572 215124 12628
rect 215852 12684 215908 12740
rect 214172 7644 214228 7700
rect 215068 7756 215124 7812
rect 211708 4172 211764 4228
rect 213164 5964 213220 6020
rect 218428 56364 218484 56420
rect 220108 59388 220164 59444
rect 221004 59388 221060 59444
rect 221788 56588 221844 56644
rect 220220 16044 220276 16100
rect 220108 14588 220164 14644
rect 216860 11340 216916 11396
rect 220108 14252 220164 14308
rect 216748 9324 216804 9380
rect 218316 10892 218372 10948
rect 215852 4956 215908 5012
rect 216972 4956 217028 5012
rect 224252 56364 224308 56420
rect 224252 29372 224308 29428
rect 225260 56364 225316 56420
rect 225148 10892 225204 10948
rect 223468 4620 223524 4676
rect 224588 7532 224644 7588
rect 222684 4508 222740 4564
rect 226492 6076 226548 6132
rect 227612 56588 227668 56644
rect 228508 7532 228564 7588
rect 229292 56476 229348 56532
rect 229292 6076 229348 6132
rect 227612 5964 227668 6020
rect 226828 4508 226884 4564
rect 228508 4396 228564 4452
rect 230300 26012 230356 26068
rect 231868 15932 231924 15988
rect 231980 16156 232036 16212
rect 230188 4396 230244 4452
rect 230300 5852 230356 5908
rect 234332 56252 234388 56308
rect 236908 56700 236964 56756
rect 238588 59388 238644 59444
rect 235340 56252 235396 56308
rect 239484 59388 239540 59444
rect 240268 55468 240324 55524
rect 238700 47852 238756 47908
rect 241948 17948 242004 18004
rect 242732 56700 242788 56756
rect 242732 17612 242788 17668
rect 238588 12684 238644 12740
rect 235228 9212 235284 9268
rect 234332 6188 234388 6244
rect 236012 7644 236068 7700
rect 233548 5852 233604 5908
rect 234108 4284 234164 4340
rect 243740 36092 243796 36148
rect 243628 7644 243684 7700
rect 243740 12572 243796 12628
rect 241724 6188 241780 6244
rect 237916 6076 237972 6132
rect 239820 4172 239876 4228
rect 246092 55468 246148 55524
rect 246092 20972 246148 21028
rect 246988 11116 247044 11172
rect 247436 11340 247492 11396
rect 245308 4284 245364 4340
rect 245532 9324 245588 9380
rect 248780 56476 248836 56532
rect 248668 2492 248724 2548
rect 248780 29372 248836 29428
rect 250348 19292 250404 19348
rect 251132 56364 251188 56420
rect 250348 16044 250404 16100
rect 252028 14364 252084 14420
rect 252140 14588 252196 14644
rect 251132 6076 251188 6132
rect 255388 56700 255444 56756
rect 253820 56364 253876 56420
rect 253708 4172 253764 4228
rect 255052 5964 255108 6020
rect 258748 56812 258804 56868
rect 257180 24332 257236 24388
rect 261212 56700 261268 56756
rect 261212 34412 261268 34468
rect 260428 6188 260484 6244
rect 260764 10892 260820 10948
rect 257068 4844 257124 4900
rect 258860 6076 258916 6132
rect 257068 4620 257124 4676
rect 262220 14252 262276 14308
rect 262108 6076 262164 6132
rect 264572 56812 264628 56868
rect 265468 44492 265524 44548
rect 266252 56476 266308 56532
rect 264572 37772 264628 37828
rect 265468 26012 265524 26068
rect 263788 4732 263844 4788
rect 264572 7532 264628 7588
rect 262668 4508 262724 4564
rect 267260 56476 267316 56532
rect 267148 16044 267204 16100
rect 267932 56252 267988 56308
rect 266252 7756 266308 7812
rect 268828 12572 268884 12628
rect 268940 15932 268996 15988
rect 267932 5964 267988 6020
rect 268380 4396 268436 4452
rect 272300 55468 272356 55524
rect 274652 55468 274708 55524
rect 274652 32732 274708 32788
rect 273868 12796 273924 12852
rect 270508 11004 270564 11060
rect 272188 5852 272244 5908
rect 272300 4620 272356 4676
rect 274092 9212 274148 9268
rect 275660 56252 275716 56308
rect 278908 54684 278964 54740
rect 279692 56476 279748 56532
rect 277228 29484 277284 29540
rect 278908 47852 278964 47908
rect 277228 17612 277284 17668
rect 275548 4508 275604 4564
rect 275996 5964 276052 6020
rect 279692 9212 279748 9268
rect 280700 29372 280756 29428
rect 280588 5964 280644 6020
rect 280700 12684 280756 12740
rect 282268 4396 282324 4452
rect 282380 20972 282436 21028
rect 285740 56700 285796 56756
rect 286412 56364 286468 56420
rect 285628 17724 285684 17780
rect 285740 17948 285796 18004
rect 283948 7532 284004 7588
rect 287308 10892 287364 10948
rect 288988 36092 289044 36148
rect 286412 7868 286468 7924
rect 287420 7644 287476 7700
rect 290668 59276 290724 59332
rect 291228 59276 291284 59332
rect 290892 56588 290948 56644
rect 290668 56476 290724 56532
rect 289100 26124 289156 26180
rect 294028 59388 294084 59444
rect 294028 56364 294084 56420
rect 294924 59388 294980 59444
rect 294252 55468 294308 55524
rect 296492 56588 296548 56644
rect 296492 27804 296548 27860
rect 298172 55468 298228 55524
rect 298172 31164 298228 31220
rect 297388 19516 297444 19572
rect 295708 17612 295764 17668
rect 297388 19292 297444 19348
rect 292348 5852 292404 5908
rect 293132 11116 293188 11172
rect 291228 4284 291284 4340
rect 296940 7756 296996 7812
rect 295036 2492 295092 2548
rect 299180 46172 299236 46228
rect 299068 12684 299124 12740
rect 300748 4284 300804 4340
rect 300860 14364 300916 14420
rect 302428 7756 302484 7812
rect 304108 59052 304164 59108
rect 302652 4172 302708 4228
rect 304780 59052 304836 59108
rect 304220 26012 304276 26068
rect 305788 15932 305844 15988
rect 305900 34412 305956 34468
rect 304108 4172 304164 4228
rect 304556 7868 304612 7924
rect 309372 55804 309428 55860
rect 309148 55468 309204 55524
rect 312508 59388 312564 59444
rect 310828 47964 310884 48020
rect 311612 55468 311668 55524
rect 307468 24556 307524 24612
rect 310828 37772 310884 37828
rect 308252 24332 308308 24388
rect 308252 4956 308308 5012
rect 310268 4956 310324 5012
rect 308364 4844 308420 4900
rect 313404 59388 313460 59444
rect 312620 55468 312676 55524
rect 312508 54572 312564 54628
rect 311612 37772 311668 37828
rect 314972 55468 315028 55524
rect 314972 36092 315028 36148
rect 314188 19292 314244 19348
rect 315980 55804 316036 55860
rect 315980 49532 316036 49588
rect 317660 56588 317716 56644
rect 317548 27692 317604 27748
rect 315868 14588 315924 14644
rect 315868 14252 315924 14308
rect 314188 6188 314244 6244
rect 319228 11116 319284 11172
rect 320908 44492 320964 44548
rect 317884 6076 317940 6132
rect 319788 4732 319844 4788
rect 321132 44492 321188 44548
rect 322700 31052 322756 31108
rect 322588 14252 322644 14308
rect 322700 16044 322756 16100
rect 325052 56700 325108 56756
rect 325948 56700 326004 56756
rect 325052 17948 325108 18004
rect 325948 12572 326004 12628
rect 324268 7644 324324 7700
rect 325500 9212 325556 9268
rect 327740 32844 327796 32900
rect 327628 12572 327684 12628
rect 330092 56700 330148 56756
rect 329308 11004 329364 11060
rect 331212 56700 331268 56756
rect 330988 55468 331044 55524
rect 333452 55468 333508 55524
rect 334348 39452 334404 39508
rect 335132 56252 335188 56308
rect 333452 37996 333508 38052
rect 332668 22764 332724 22820
rect 332780 32732 332836 32788
rect 330092 9324 330148 9380
rect 329420 6188 329476 6244
rect 331212 4620 331268 4676
rect 334348 12796 334404 12852
rect 336140 56252 336196 56308
rect 337708 12796 337764 12852
rect 336028 11004 336084 11060
rect 335132 5740 335188 5796
rect 338828 5740 338884 5796
rect 336924 4508 336980 4564
rect 341068 59388 341124 59444
rect 339388 2604 339444 2660
rect 339500 29484 339556 29540
rect 341740 59388 341796 59444
rect 341180 21084 341236 21140
rect 342748 54684 342804 54740
rect 341068 6076 341124 6132
rect 344428 56812 344484 56868
rect 342860 46396 342916 46452
rect 347788 54908 347844 54964
rect 349468 59388 349524 59444
rect 346220 44716 346276 44772
rect 346108 34524 346164 34580
rect 346108 29372 346164 29428
rect 344540 5964 344596 6020
rect 350364 59388 350420 59444
rect 349580 53116 349636 53172
rect 351148 29484 351204 29540
rect 351932 56700 351988 56756
rect 354620 58044 354676 58100
rect 354508 36204 354564 36260
rect 355292 56812 355348 56868
rect 352828 19404 352884 19460
rect 351932 17836 351988 17892
rect 352828 17948 352884 18004
rect 349468 16044 349524 16100
rect 351148 17724 351204 17780
rect 350252 7532 350308 7588
rect 348348 4396 348404 4452
rect 356188 48076 356244 48132
rect 356972 56476 357028 56532
rect 355292 17724 355348 17780
rect 355964 10892 356020 10948
rect 357868 41356 357924 41412
rect 359660 51436 359716 51492
rect 359548 39564 359604 39620
rect 359548 27804 359604 27860
rect 356972 8092 357028 8148
rect 357868 26124 357924 26180
rect 361228 20972 361284 21028
rect 362012 56364 362068 56420
rect 361676 8092 361732 8148
rect 362908 56364 362964 56420
rect 362012 6300 362068 6356
rect 366268 56812 366324 56868
rect 364700 56476 364756 56532
rect 365596 56364 365652 56420
rect 365596 51324 365652 51380
rect 364588 5964 364644 6020
rect 364700 31164 364756 31220
rect 363580 5852 363636 5908
rect 368060 46284 368116 46340
rect 369628 29372 369684 29428
rect 370412 56588 370468 56644
rect 367948 26124 368004 26180
rect 367948 17612 368004 17668
rect 367388 6300 367444 6356
rect 372092 56812 372148 56868
rect 372092 42924 372148 42980
rect 371308 31164 371364 31220
rect 370412 7868 370468 7924
rect 371308 19516 371364 19572
rect 373100 53004 373156 53060
rect 374668 34412 374724 34468
rect 374780 46172 374836 46228
rect 372988 7532 373044 7588
rect 374668 12684 374724 12740
rect 373324 4956 373380 5012
rect 374780 4956 374836 5012
rect 378140 57932 378196 57988
rect 381388 55468 381444 55524
rect 379708 22652 379764 22708
rect 379820 26012 379876 26068
rect 378028 9212 378084 9268
rect 378812 7756 378868 7812
rect 376348 2492 376404 2548
rect 376908 4284 376964 4340
rect 384748 56700 384804 56756
rect 386428 59388 386484 59444
rect 383180 56588 383236 56644
rect 383852 55468 383908 55524
rect 383852 46172 383908 46228
rect 383068 24444 383124 24500
rect 387324 59388 387380 59444
rect 386540 56364 386596 56420
rect 388332 37884 388388 37940
rect 389788 49532 389844 49588
rect 388108 37772 388164 37828
rect 386428 24332 386484 24388
rect 386540 24556 386596 24612
rect 383068 15932 383124 15988
rect 382620 4172 382676 4228
rect 390348 56700 390404 56756
rect 390348 49644 390404 49700
rect 389900 47852 389956 47908
rect 393148 56700 393204 56756
rect 391580 55468 391636 55524
rect 393596 56588 393652 56644
rect 391468 10892 391524 10948
rect 391580 47964 391636 48020
rect 393596 47964 393652 48020
rect 393932 55468 393988 55524
rect 393932 44604 393988 44660
rect 394828 54572 394884 54628
rect 393148 36092 393204 36148
rect 394940 32732 394996 32788
rect 398188 56588 398244 56644
rect 396620 51212 396676 51268
rect 396508 17612 396564 17668
rect 396620 19292 396676 19348
rect 401660 55468 401716 55524
rect 403228 49532 403284 49588
rect 401548 37772 401604 37828
rect 403228 27692 403284 27748
rect 399868 14364 399924 14420
rect 399980 14588 400036 14644
rect 401660 7868 401716 7924
rect 405020 19292 405076 19348
rect 406588 44492 406644 44548
rect 404908 4732 404964 4788
rect 405468 11116 405524 11172
rect 407372 55468 407428 55524
rect 407372 44492 407428 44548
rect 406700 27804 406756 27860
rect 408268 4620 408324 4676
rect 408380 31052 408436 31108
rect 410060 54796 410116 54852
rect 409948 5852 410004 5908
rect 410060 14252 410116 14308
rect 412412 56700 412468 56756
rect 413308 15932 413364 15988
rect 416668 54684 416724 54740
rect 415100 41244 415156 41300
rect 418348 26012 418404 26068
rect 418460 32844 418516 32900
rect 414988 12684 415044 12740
rect 415772 12572 415828 12628
rect 414988 9324 415044 9380
rect 412412 7644 412468 7700
rect 413084 7756 413140 7812
rect 411628 4508 411684 4564
rect 415772 4956 415828 5012
rect 416892 4956 416948 5012
rect 420140 54572 420196 54628
rect 421708 37996 421764 38052
rect 420028 4396 420084 4452
rect 420700 6188 420756 6244
rect 421820 36092 421876 36148
rect 423500 52892 423556 52948
rect 426748 56812 426804 56868
rect 425068 27692 425124 27748
rect 427532 56252 427588 56308
rect 425068 22764 425124 22820
rect 423388 4284 423444 4340
rect 423500 17836 423556 17892
rect 428428 56252 428484 56308
rect 427532 6748 427588 6804
rect 428428 39452 428484 39508
rect 428540 31052 428596 31108
rect 431788 56700 431844 56756
rect 433468 59388 433524 59444
rect 432572 56476 432628 56532
rect 432572 17836 432628 17892
rect 430108 12572 430164 12628
rect 432124 11004 432180 11060
rect 430220 6748 430276 6804
rect 434140 59388 434196 59444
rect 441868 438620 441924 438676
rect 440188 41132 440244 41188
rect 440300 46396 440356 46452
rect 436828 21868 436884 21924
rect 433580 14252 433636 14308
rect 436828 21084 436884 21140
rect 433468 4172 433524 4228
rect 433580 12796 433636 12852
rect 435932 2604 435988 2660
rect 439740 6076 439796 6132
rect 442652 430108 442708 430164
rect 444332 231868 444388 231924
rect 446012 440524 446068 440580
rect 474348 590492 474404 590548
rect 518476 593180 518532 593236
rect 540540 593068 540596 593124
rect 495628 461244 495684 461300
rect 454412 457772 454468 457828
rect 486332 455532 486388 455588
rect 484652 455420 484708 455476
rect 481292 455308 481348 455364
rect 477932 453740 477988 453796
rect 476252 452060 476308 452116
rect 466172 450716 466228 450772
rect 464492 450492 464548 450548
rect 459452 450268 459508 450324
rect 456092 445452 456148 445508
rect 451052 443772 451108 443828
rect 449372 441980 449428 442036
rect 449372 416668 449428 416724
rect 451052 362908 451108 362964
rect 454412 441868 454468 441924
rect 447692 270508 447748 270564
rect 446012 204988 446068 205044
rect 454412 178108 454468 178164
rect 467852 445564 467908 445620
rect 467852 389788 467908 389844
rect 466172 349468 466228 349524
rect 464492 310828 464548 310884
rect 459452 218428 459508 218484
rect 456092 112588 456148 112644
rect 479612 447244 479668 447300
rect 487788 455308 487844 455364
rect 487788 454412 487844 454468
rect 486332 376348 486388 376404
rect 496412 447020 496468 447076
rect 484652 336028 484708 336084
rect 481292 297388 481348 297444
rect 479612 257068 479668 257124
rect 477932 137788 477988 137844
rect 476252 99148 476308 99204
rect 584892 590492 584948 590548
rect 593292 590492 593348 590548
rect 593068 562156 593124 562212
rect 593180 522508 593236 522564
rect 593292 467852 593348 467908
rect 593740 473788 593796 473844
rect 593180 466172 593236 466228
rect 593404 467068 593460 467124
rect 593068 464492 593124 464548
rect 593180 465388 593236 465444
rect 590492 448588 590548 448644
rect 588812 446908 588868 446964
rect 588812 443436 588868 443492
rect 561148 442652 561204 442708
rect 593068 440188 593124 440244
rect 593068 403788 593124 403844
rect 590492 192332 590548 192388
rect 496412 58828 496468 58884
rect 458668 58044 458724 58100
rect 446012 56812 446068 56868
rect 444332 56588 444388 56644
rect 441868 8428 441924 8484
rect 443548 17724 443604 17780
rect 454412 56700 454468 56756
rect 448588 54908 448644 54964
rect 446012 39452 446068 39508
rect 446908 44716 446964 44772
rect 445228 34524 445284 34580
rect 444332 9324 444388 9380
rect 450268 53116 450324 53172
rect 454412 32844 454468 32900
rect 453628 29484 453684 29540
rect 451948 16044 452004 16100
rect 456092 19404 456148 19460
rect 493948 57932 494004 57988
rect 484652 56364 484708 56420
rect 465388 51436 465444 51492
rect 462028 48076 462084 48132
rect 460348 36204 460404 36260
rect 456092 4956 456148 5012
rect 456988 4956 457044 5012
rect 463708 41356 463764 41412
rect 472108 51324 472164 51380
rect 467068 39564 467124 39620
rect 468748 20972 468804 21028
rect 480508 46284 480564 46340
rect 477148 42924 477204 42980
rect 475468 17836 475524 17892
rect 474012 5964 474068 6020
rect 478828 26124 478884 26180
rect 482188 29372 482244 29428
rect 487228 53004 487284 53060
rect 484652 5964 484708 6020
rect 485548 31164 485604 31220
rect 490588 34412 490644 34468
rect 489244 7532 489300 7588
rect 493052 2492 493108 2548
rect 570332 56252 570388 56308
rect 544348 54796 544404 54852
rect 522508 51212 522564 51268
rect 505708 49644 505764 49700
rect 502348 47964 502404 48020
rect 500668 46172 500724 46228
rect 497308 22652 497364 22708
rect 496860 9212 496916 9268
rect 504028 24444 504084 24500
rect 514108 47852 514164 47908
rect 512428 37884 512484 37940
rect 509068 24332 509124 24388
rect 508284 5964 508340 6020
rect 515788 44604 515844 44660
rect 520828 32732 520884 32788
rect 517804 10892 517860 10948
rect 519708 7644 519764 7700
rect 534268 49532 534324 49588
rect 530908 44492 530964 44548
rect 523292 17612 523348 17668
rect 529228 14364 529284 14420
rect 527324 9324 527380 9380
rect 523292 4956 523348 5012
rect 525420 4956 525476 5012
rect 532588 37772 532644 37828
rect 539308 27804 539364 27860
rect 537628 19292 537684 19348
rect 536844 4732 536900 4788
rect 554428 54684 554484 54740
rect 551068 41244 551124 41300
rect 549388 15932 549444 15988
rect 542668 4620 542724 4676
rect 546364 5852 546420 5908
rect 548268 4508 548324 4564
rect 552748 12684 552804 12740
rect 560252 54572 560308 54628
rect 557788 26012 557844 26068
rect 566188 52892 566244 52948
rect 562828 36092 562884 36148
rect 560252 4956 560308 5012
rect 561596 4956 561652 5012
rect 559692 4396 559748 4452
rect 565404 4284 565460 4340
rect 567868 27692 567924 27748
rect 590492 42812 590548 42868
rect 570332 10108 570388 10164
rect 571228 39452 571284 39508
rect 579628 32844 579684 32900
rect 574588 31052 574644 31108
rect 573020 10108 573076 10164
rect 576268 12572 576324 12628
rect 593292 445228 593348 445284
rect 593628 458668 593684 458724
rect 593516 456988 593572 457044
rect 594076 470428 594132 470484
rect 593852 462028 593908 462084
rect 593964 451948 594020 452004
rect 594188 460348 594244 460404
rect 594188 324492 594244 324548
rect 594300 443548 594356 443604
rect 594076 284844 594132 284900
rect 593964 245196 594020 245252
rect 593852 165900 593908 165956
rect 593740 152684 593796 152740
rect 593628 126252 593684 126308
rect 593516 86604 593572 86660
rect 593404 73388 593460 73444
rect 593292 46956 593348 47012
rect 593180 33740 593236 33796
rect 590492 20524 590548 20580
rect 581308 14252 581364 14308
rect 594300 7308 594356 7364
rect 584444 4172 584500 4228
<< metal3 >>
rect 231858 593404 231868 593460
rect 231924 593404 451612 593460
rect 451668 593404 451678 593460
rect 55346 593292 55356 593348
rect 55412 593292 288988 593348
rect 289044 593292 289054 593348
rect 224242 593180 224252 593236
rect 224308 593180 518476 593236
rect 518532 593180 518542 593236
rect 215058 593068 215068 593124
rect 215124 593068 540540 593124
rect 540596 593068 540606 593124
rect 99474 591276 99484 591332
rect 99540 591276 104972 591332
rect 105028 591276 105038 591332
rect 427522 590828 427532 590884
rect 427588 590828 430220 590884
rect 430276 590828 430286 590884
rect 187730 590604 187740 590660
rect 187796 590604 188972 590660
rect 189028 590604 189038 590660
rect 242722 590604 242732 590660
rect 242788 590604 386092 590660
rect 386148 590604 386158 590660
rect 33282 590492 33292 590548
rect 33348 590492 274652 590548
rect 274708 590492 274718 590548
rect 303202 590492 303212 590548
rect 303268 590492 364028 590548
rect 364084 590492 364094 590548
rect 454402 590492 454412 590548
rect 454468 590492 474348 590548
rect 474404 590492 474414 590548
rect 584882 590492 584892 590548
rect 584948 590492 593292 590548
rect 593348 590492 593358 590548
rect 595560 588644 597000 588840
rect 595420 588616 597000 588644
rect 595420 588588 595672 588616
rect 595420 588532 595476 588588
rect 595420 588476 595700 588532
rect 595644 588084 595700 588476
rect 207442 588028 207452 588084
rect 207508 588028 595700 588084
rect -960 587188 480 587384
rect -960 587160 532 587188
rect 392 587132 532 587160
rect 476 587076 532 587132
rect 364 587020 532 587076
rect 364 586404 420 587020
rect 364 586348 299068 586404
rect 299124 586348 299134 586404
rect 595560 575428 597000 575624
rect 208562 575372 208572 575428
rect 208628 575372 263788 575428
rect 263844 575372 263854 575428
rect 595420 575400 597000 575428
rect 595420 575372 595672 575400
rect 595420 575316 595476 575372
rect 595420 575260 595700 575316
rect 595644 574644 595700 575260
rect 208338 574588 208348 574644
rect 208404 574588 595700 574644
rect -960 573076 480 573272
rect -960 573048 11788 573076
rect 392 573020 11788 573048
rect 11732 572964 11788 573020
rect 11732 572908 305788 572964
rect 305844 572908 305864 572964
rect 595560 562212 597000 562408
rect 593058 562156 593068 562212
rect 593124 562184 597000 562212
rect 593124 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 532 558964
rect 392 558908 532 558936
rect 476 558852 532 558908
rect 364 558796 532 558852
rect 364 557844 420 558796
rect 364 557788 12572 557844
rect 12628 557788 12638 557844
rect 595560 548996 597000 549192
rect 595420 548968 597000 548996
rect 595420 548940 595672 548968
rect 595420 548884 595476 548940
rect 595420 548828 595700 548884
rect 595644 547764 595700 548828
rect 194898 547708 194908 547764
rect 194964 547708 595700 547764
rect -960 544852 480 545048
rect -960 544824 532 544852
rect 392 544796 532 544824
rect 476 544740 532 544796
rect 364 544684 532 544740
rect 364 544404 420 544684
rect 364 544348 308252 544404
rect 308308 544348 308318 544404
rect 595560 535780 597000 535976
rect 595420 535752 597000 535780
rect 595420 535724 595672 535752
rect 595420 535668 595476 535724
rect 595420 535612 595700 535668
rect 595644 534324 595700 535612
rect 198258 534268 198268 534324
rect 198324 534268 595700 534324
rect -960 530740 480 530936
rect -960 530712 5852 530740
rect 392 530684 5852 530712
rect 5908 530684 5918 530740
rect 595560 522564 597000 522760
rect 593170 522508 593180 522564
rect 593236 522536 597000 522564
rect 593236 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 4172 516628
rect 392 516572 4172 516600
rect 4228 516572 4238 516628
rect 595560 509348 597000 509544
rect 587972 509320 597000 509348
rect 587972 509292 595672 509320
rect 587972 509124 588028 509292
rect 194002 509068 194012 509124
rect 194068 509068 588028 509124
rect 250338 503132 250348 503188
rect 250404 503132 319228 503188
rect 319284 503132 319294 503188
rect -960 502516 480 502712
rect -960 502488 11788 502516
rect 392 502460 11788 502488
rect 11732 502404 11788 502460
rect 11732 502348 212492 502404
rect 212548 502348 212558 502404
rect 595560 496132 597000 496328
rect 595420 496104 597000 496132
rect 595420 496076 595672 496104
rect 595420 496020 595476 496076
rect 595420 495964 595700 496020
rect 595644 495684 595700 495964
rect 189858 495628 189868 495684
rect 189924 495628 595700 495684
rect -960 488404 480 488600
rect -960 488376 532 488404
rect 392 488348 532 488376
rect 476 488292 532 488348
rect 364 488236 532 488292
rect 364 487284 420 488236
rect 364 487228 325052 487284
rect 325108 487228 325118 487284
rect 595560 482916 597000 483112
rect 595420 482888 597000 482916
rect 595420 482860 595672 482888
rect 595420 482804 595476 482860
rect 595420 482748 595700 482804
rect 595644 482244 595700 482748
rect 185602 482188 185612 482244
rect 185668 482188 595700 482244
rect 212482 476252 212492 476308
rect 212548 476252 319228 476308
rect 319284 476252 319294 476308
rect 120978 474572 120988 474628
rect 121044 474572 280588 474628
rect 280644 474572 280654 474628
rect -960 474292 480 474488
rect -960 474264 532 474292
rect 392 474236 532 474264
rect 476 474180 532 474236
rect 364 474124 532 474180
rect 364 473844 420 474124
rect 364 473788 14252 473844
rect 14308 473788 14318 473844
rect 97458 473788 97468 473844
rect 97524 473788 593740 473844
rect 593796 473788 593806 473844
rect 188962 472892 188972 472948
rect 189028 472892 270508 472948
rect 270564 472892 270574 472948
rect 17602 472108 17612 472164
rect 17668 472108 409948 472164
rect 410004 472108 410014 472164
rect 253698 471212 253708 471268
rect 253764 471212 260428 471268
rect 260484 471212 260494 471268
rect 22642 470540 22652 470596
rect 22708 470540 393148 470596
rect 393204 470540 393214 470596
rect 134418 470428 134428 470484
rect 134484 470428 594076 470484
rect 594132 470428 594142 470484
rect 595560 469700 597000 469896
rect 595420 469672 597000 469700
rect 595420 469644 595672 469672
rect 595420 469588 595476 469644
rect 238578 469532 238588 469588
rect 238644 469532 427532 469588
rect 427588 469532 427598 469588
rect 595420 469532 595700 469588
rect 2482 468860 2492 468916
rect 2548 468860 413308 468916
rect 413364 468860 413374 468916
rect 595644 468804 595700 469532
rect 176418 468748 176428 468804
rect 176484 468748 595700 468804
rect 211698 467852 211708 467908
rect 211764 467852 593292 467908
rect 593348 467852 593358 467908
rect 27682 467180 27692 467236
rect 27748 467180 403228 467236
rect 403284 467180 403294 467236
rect 78978 467068 78988 467124
rect 79044 467068 593404 467124
rect 593460 467068 593470 467124
rect 191538 466172 191548 466228
rect 191604 466172 593180 466228
rect 593236 466172 593246 466228
rect 19282 465500 19292 465556
rect 19348 465500 364588 465556
rect 364644 465500 364654 465556
rect 68898 465388 68908 465444
rect 68964 465388 593180 465444
rect 593236 465388 593246 465444
rect 230178 464604 230188 464660
rect 230244 464604 267148 464660
rect 267204 464604 267214 464660
rect 201618 464492 201628 464548
rect 201684 464492 593068 464548
rect 593124 464492 593134 464548
rect 36082 463820 36092 463876
rect 36148 463820 371308 463876
rect 371364 463820 371374 463876
rect 9202 463708 9212 463764
rect 9268 463708 406588 463764
rect 406644 463708 406654 463764
rect 257058 463036 257068 463092
rect 257124 463036 297388 463092
rect 297444 463036 297454 463092
rect 246978 462924 246988 462980
rect 247044 462924 303212 462980
rect 303268 462924 303278 462980
rect 5842 462812 5852 462868
rect 5908 462812 315868 462868
rect 315924 462812 315934 462868
rect 127698 462140 127708 462196
rect 127764 462140 447692 462196
rect 447748 462140 447758 462196
rect 104178 462028 104188 462084
rect 104244 462028 593852 462084
rect 593908 462028 593918 462084
rect 104962 461356 104972 461412
rect 105028 461356 287308 461412
rect 287364 461356 287374 461412
rect 228498 461244 228508 461300
rect 228564 461244 495628 461300
rect 495684 461244 495694 461300
rect 14242 461132 14252 461188
rect 14308 461132 322588 461188
rect 322644 461132 322654 461188
rect -960 460180 480 460376
rect 142930 460348 142940 460404
rect 142996 460348 594188 460404
rect 594244 460348 594254 460404
rect -960 460152 532 460180
rect 392 460124 532 460152
rect 476 460068 532 460124
rect 364 460012 532 460068
rect 364 458836 420 460012
rect 253698 459676 253708 459732
rect 253764 459676 275548 459732
rect 275604 459676 275614 459732
rect 243618 459564 243628 459620
rect 243684 459564 341068 459620
rect 341124 459564 341134 459620
rect 12562 459452 12572 459508
rect 12628 459452 302428 459508
rect 302484 459452 302494 459508
rect 117618 458892 117628 458948
rect 117684 458892 444332 458948
rect 444388 458892 444398 458948
rect 364 458780 246092 458836
rect 246148 458780 246158 458836
rect 94098 458668 94108 458724
rect 94164 458668 593628 458724
rect 593684 458668 593694 458724
rect 142818 457996 142828 458052
rect 142884 457996 273868 458052
rect 273924 457996 273934 458052
rect 274642 457996 274652 458052
rect 274708 457996 295708 458052
rect 295764 457996 295774 458052
rect 235218 457884 235228 457940
rect 235284 457884 408268 457940
rect 408324 457884 408334 457940
rect 225138 457772 225148 457828
rect 225204 457772 454412 457828
rect 454468 457772 454478 457828
rect 15922 457100 15932 457156
rect 15988 457100 361228 457156
rect 361284 457100 361294 457156
rect 85698 456988 85708 457044
rect 85764 456988 593516 457044
rect 593572 456988 593582 457044
rect 595560 456484 597000 456680
rect 595420 456456 597000 456484
rect 595420 456428 595672 456456
rect 595420 456372 595476 456428
rect 595420 456316 595700 456372
rect 14242 455644 14252 455700
rect 14308 455644 332668 455700
rect 332724 455644 332734 455700
rect 159618 455532 159628 455588
rect 159684 455532 486332 455588
rect 486388 455532 486398 455588
rect 149538 455420 149548 455476
rect 149604 455420 484652 455476
rect 484708 455420 484718 455476
rect 595644 455364 595700 456316
rect 141138 455308 141148 455364
rect 141204 455308 481292 455364
rect 481348 455308 481358 455364
rect 487778 455308 487788 455364
rect 487844 455308 595700 455364
rect 246082 454524 246092 454580
rect 246148 454524 329308 454580
rect 329364 454524 329384 454580
rect 179778 454412 179788 454468
rect 179844 454412 487788 454468
rect 487844 454412 487854 454468
rect 52882 453852 52892 453908
rect 52948 453852 386428 453908
rect 386484 453852 386494 453908
rect 100818 453740 100828 453796
rect 100884 453740 477932 453796
rect 477988 453740 477998 453796
rect 44482 453628 44492 453684
rect 44548 453628 423388 453684
rect 423444 453628 423464 453684
rect 31042 452284 31052 452340
rect 31108 452284 354508 452340
rect 354564 452284 354574 452340
rect 41122 452172 41132 452228
rect 41188 452172 384748 452228
rect 384804 452172 384814 452228
rect 92418 452060 92428 452116
rect 92484 452060 476252 452116
rect 476308 452060 476318 452116
rect 124338 451948 124348 452004
rect 124404 451948 593964 452004
rect 594020 451948 594030 452004
rect 146178 450716 146188 450772
rect 146244 450716 466172 450772
rect 466228 450716 466238 450772
rect 54562 450604 54572 450660
rect 54628 450604 378028 450660
rect 378084 450604 378094 450660
rect 137778 450492 137788 450548
rect 137844 450492 464492 450548
rect 464548 450492 464558 450548
rect 37762 450380 37772 450436
rect 37828 450380 374668 450436
rect 374724 450380 374734 450436
rect 120978 450268 120988 450324
rect 121044 450268 459452 450324
rect 459508 450268 459518 450324
rect 44594 449036 44604 449092
rect 44660 449036 344428 449092
rect 344484 449036 344494 449092
rect 51202 448924 51212 448980
rect 51268 448924 396508 448980
rect 396564 448924 396574 448980
rect 29362 448812 29372 448868
rect 29428 448812 389788 448868
rect 389844 448812 389854 448868
rect 32722 448700 32732 448756
rect 32788 448700 399868 448756
rect 399924 448700 399944 448756
rect 170482 448588 170492 448644
rect 170548 448588 590492 448644
rect 590548 448588 590558 448644
rect 325042 448476 325052 448532
rect 325108 448476 325948 448532
rect 326004 448476 326014 448532
rect 46162 447356 46172 447412
rect 46228 447356 351148 447412
rect 351204 447356 351214 447412
rect 131058 447244 131068 447300
rect 131124 447244 479612 447300
rect 479668 447244 479678 447300
rect 5842 447132 5852 447188
rect 5908 447132 367948 447188
rect 368004 447132 368014 447188
rect 82338 447020 82348 447076
rect 82404 447020 496412 447076
rect 496468 447020 496478 447076
rect 173058 446908 173068 446964
rect 173124 446908 588812 446964
rect 588868 446908 588878 446964
rect -960 446068 480 446264
rect -960 446040 532 446068
rect 392 446012 532 446040
rect 476 445956 532 446012
rect 364 445900 532 445956
rect 364 445396 420 445900
rect 47842 445676 47852 445732
rect 47908 445676 342524 445732
rect 342580 445676 342590 445732
rect 157378 445564 157388 445620
rect 157444 445564 467852 445620
rect 467908 445564 467918 445620
rect 89170 445452 89180 445508
rect 89236 445452 456092 445508
rect 456148 445452 456158 445508
rect 364 445340 336028 445396
rect 336084 445340 336094 445396
rect 76178 445228 76188 445284
rect 76244 445228 593292 445284
rect 593348 445228 593358 445284
rect 186610 444332 186620 444388
rect 186676 444332 194012 444388
rect 194068 444332 194078 444388
rect 183362 444108 183372 444164
rect 183428 444108 185612 444164
rect 185668 444108 185678 444164
rect 206098 444108 206108 444164
rect 206164 444108 207452 444164
rect 207508 444108 207518 444164
rect 241826 444108 241836 444164
rect 241892 444108 242732 444164
rect 242788 444108 242798 444164
rect 167122 443996 167132 444052
rect 167188 443996 442652 444052
rect 442708 443996 442718 444052
rect 56242 443884 56252 443940
rect 56308 443884 349020 443940
rect 349076 443884 349086 443940
rect 154130 443772 154140 443828
rect 154196 443772 451052 443828
rect 451108 443772 451118 443828
rect 12562 443660 12572 443716
rect 12628 443660 358764 443716
rect 358820 443660 358830 443716
rect 66434 443548 66444 443604
rect 66500 443548 594300 443604
rect 594356 443548 594366 443604
rect 588802 443436 588812 443492
rect 588868 443464 595672 443492
rect 588868 443436 597000 443464
rect 222338 443212 222348 443268
rect 222404 443212 224252 443268
rect 224308 443212 224318 443268
rect 595560 443240 597000 443436
rect 164658 443100 164668 443156
rect 164724 443100 277564 443156
rect 277620 443100 277630 443156
rect 308242 443100 308252 443156
rect 308308 443100 310044 443156
rect 310100 443100 310110 443156
rect 77298 442988 77308 443044
rect 77364 442988 284060 443044
rect 284116 442988 284126 443044
rect 10098 442876 10108 442932
rect 10164 442876 293804 442932
rect 293860 442876 293870 442932
rect 4162 442764 4172 442820
rect 4228 442764 313292 442820
rect 313348 442764 313358 442820
rect 108658 442652 108668 442708
rect 108724 442652 170492 442708
rect 170548 442652 170558 442708
rect 219090 442652 219100 442708
rect 219156 442652 561148 442708
rect 561204 442652 561214 442708
rect 426962 442092 426972 442148
rect 427028 442092 440188 442148
rect 440244 442092 440254 442148
rect 170370 441980 170380 442036
rect 170436 441980 449372 442036
rect 449428 441980 449438 442036
rect 60386 441868 60396 441924
rect 60452 441868 72940 441924
rect 72996 441868 73006 441924
rect 111906 441868 111916 441924
rect 111972 441868 454412 441924
rect 454468 441868 454478 441924
rect 59602 440636 59612 440692
rect 59668 440636 339276 440692
rect 339332 440636 339342 440692
rect 115154 440524 115164 440580
rect 115220 440524 446012 440580
rect 446068 440524 446078 440580
rect 49522 440412 49532 440468
rect 49588 440412 417228 440468
rect 417284 440412 417294 440468
rect 34402 440300 34412 440356
rect 34468 440300 420476 440356
rect 420532 440300 420542 440356
rect 163874 440188 163884 440244
rect 163940 440188 593068 440244
rect 593124 440188 593134 440244
rect 376292 439292 381500 439348
rect 381556 439292 381566 439348
rect 430210 439292 430220 439348
rect 430276 439292 430286 439348
rect 433430 439292 433468 439348
rect 433524 439292 433534 439348
rect 376292 438564 376348 439292
rect 430220 438676 430276 439292
rect 430220 438620 441868 438676
rect 441924 438620 441934 438676
rect 10882 438508 10892 438564
rect 10948 438508 376348 438564
rect 433458 438508 433468 438564
rect 433524 438508 436828 438564
rect 436884 438508 436894 438564
rect -960 431956 480 432152
rect -960 431928 11788 431956
rect 392 431900 11788 431928
rect 11732 431844 11788 431900
rect 11732 431788 14252 431844
rect 14308 431788 14318 431844
rect 595560 430164 597000 430248
rect 442642 430108 442652 430164
rect 442708 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 532 417844
rect 392 417788 532 417816
rect 476 417732 532 417788
rect 364 417676 532 417732
rect 364 416724 420 417676
rect 595560 416836 597000 417032
rect 587972 416808 597000 416836
rect 587972 416780 595672 416808
rect 587972 416724 588028 416780
rect 364 416668 59612 416724
rect 59668 416668 59678 416724
rect 449362 416668 449372 416724
rect 449428 416668 588028 416724
rect -960 403732 480 403928
rect 593058 403788 593068 403844
rect 593124 403816 595672 403844
rect 593124 403788 597000 403816
rect -960 403704 532 403732
rect 392 403676 532 403704
rect 476 403620 532 403676
rect 364 403564 532 403620
rect 595560 403592 597000 403788
rect 364 403284 420 403564
rect 364 403228 44604 403284
rect 44660 403228 44670 403284
rect 595560 390404 597000 390600
rect 595420 390376 597000 390404
rect 595420 390348 595672 390376
rect 595420 390292 595476 390348
rect 595420 390236 595700 390292
rect 595644 389844 595700 390236
rect -960 389620 480 389816
rect 467842 389788 467852 389844
rect 467908 389788 595700 389844
rect -960 389592 532 389620
rect 392 389564 532 389592
rect 476 389508 532 389564
rect 364 389452 532 389508
rect 364 388164 420 389452
rect 364 388108 47852 388164
rect 47908 388108 47918 388164
rect 595560 377188 597000 377384
rect 595420 377160 597000 377188
rect 595420 377132 595672 377160
rect 595420 377076 595476 377132
rect 595420 377020 595700 377076
rect 595644 376404 595700 377020
rect 486322 376348 486332 376404
rect 486388 376348 595700 376404
rect -960 375508 480 375704
rect -960 375480 532 375508
rect 392 375452 532 375480
rect 476 375396 532 375452
rect 364 375340 532 375396
rect 364 374724 420 375340
rect 364 374668 56252 374724
rect 56308 374668 56318 374724
rect 595560 363972 597000 364168
rect 595420 363944 597000 363972
rect 595420 363916 595672 363944
rect 595420 363860 595476 363916
rect 595420 363804 595700 363860
rect 595644 362964 595700 363804
rect 451042 362908 451052 362964
rect 451108 362908 595700 362964
rect -960 361396 480 361592
rect -960 361368 11788 361396
rect 392 361340 11788 361368
rect 11732 361284 11788 361340
rect 11732 361228 31052 361284
rect 31108 361228 31118 361284
rect 595560 350756 597000 350952
rect 595420 350728 597000 350756
rect 595420 350700 595672 350728
rect 595420 350644 595476 350700
rect 595420 350588 595700 350644
rect 595644 349524 595700 350588
rect 466162 349468 466172 349524
rect 466228 349468 595700 349524
rect -960 347284 480 347480
rect -960 347256 532 347284
rect 392 347228 532 347256
rect 476 347172 532 347228
rect 364 347116 532 347172
rect 364 346164 420 347116
rect 364 346108 46172 346164
rect 46228 346108 46238 346164
rect 595560 337540 597000 337736
rect 595420 337512 597000 337540
rect 595420 337484 595672 337512
rect 595420 337428 595476 337484
rect 595420 337372 595700 337428
rect 595644 336084 595700 337372
rect 484642 336028 484652 336084
rect 484708 336028 595700 336084
rect -960 333172 480 333368
rect -960 333144 532 333172
rect 392 333116 532 333144
rect 476 333060 532 333116
rect 364 333004 532 333060
rect 364 332724 420 333004
rect 364 332668 12572 332724
rect 12628 332668 12638 332724
rect 594178 324492 594188 324548
rect 594244 324520 595672 324548
rect 594244 324492 597000 324520
rect 595560 324296 597000 324492
rect -960 319060 480 319256
rect -960 319032 532 319060
rect 392 319004 532 319032
rect 476 318948 532 319004
rect 364 318892 532 318948
rect 364 317604 420 318892
rect 364 317548 19292 317604
rect 19348 317548 19358 317604
rect 595560 311108 597000 311304
rect 587972 311080 597000 311108
rect 587972 311052 595672 311080
rect 587972 310884 588028 311052
rect 464482 310828 464492 310884
rect 464548 310828 588028 310884
rect -960 304948 480 305144
rect -960 304920 532 304948
rect 392 304892 532 304920
rect 476 304836 532 304892
rect 364 304780 532 304836
rect 364 304164 420 304780
rect 364 304108 15932 304164
rect 15988 304108 15998 304164
rect 595560 297892 597000 298088
rect 595420 297864 597000 297892
rect 595420 297836 595672 297864
rect 595420 297780 595476 297836
rect 595420 297724 595700 297780
rect 595644 297444 595700 297724
rect 481282 297388 481292 297444
rect 481348 297388 595700 297444
rect 392 291032 5852 291060
rect -960 291004 5852 291032
rect 5908 291004 5918 291060
rect -960 290808 480 291004
rect 594066 284844 594076 284900
rect 594132 284872 595672 284900
rect 594132 284844 597000 284872
rect 595560 284648 597000 284844
rect -960 276724 480 276920
rect -960 276696 532 276724
rect 392 276668 532 276696
rect 476 276612 532 276668
rect 364 276556 532 276612
rect 364 275604 420 276556
rect 364 275548 37772 275604
rect 37828 275548 37838 275604
rect 595560 271460 597000 271656
rect 595420 271432 597000 271460
rect 595420 271404 595672 271432
rect 595420 271348 595476 271404
rect 595420 271292 595700 271348
rect 595644 270564 595700 271292
rect 447682 270508 447692 270564
rect 447748 270508 595700 270564
rect -960 262612 480 262808
rect -960 262584 532 262612
rect 392 262556 532 262584
rect 476 262500 532 262556
rect 364 262444 532 262500
rect 364 262164 420 262444
rect 364 262108 36092 262164
rect 36148 262108 36158 262164
rect 595560 258244 597000 258440
rect 595420 258216 597000 258244
rect 595420 258188 595672 258216
rect 595420 258132 595476 258188
rect 595420 258076 595700 258132
rect 595644 257124 595700 258076
rect 479602 257068 479612 257124
rect 479668 257068 595700 257124
rect -960 248500 480 248696
rect -960 248472 532 248500
rect 392 248444 532 248472
rect 476 248388 532 248444
rect 364 248332 532 248388
rect 364 247044 420 248332
rect 364 246988 54572 247044
rect 54628 246988 54638 247044
rect 593954 245196 593964 245252
rect 594020 245224 595672 245252
rect 594020 245196 597000 245224
rect 595560 245000 597000 245196
rect -960 234388 480 234584
rect -960 234360 532 234388
rect 392 234332 532 234360
rect 476 234276 532 234332
rect 364 234220 532 234276
rect 364 233604 420 234220
rect 364 233548 41132 233604
rect 41188 233548 41198 233604
rect 595560 231924 597000 232008
rect 444322 231868 444332 231924
rect 444388 231868 597000 231924
rect 595560 231784 597000 231868
rect 392 220472 10892 220500
rect -960 220444 10892 220472
rect 10948 220444 10958 220500
rect -960 220248 480 220444
rect 595560 218596 597000 218792
rect 587972 218568 597000 218596
rect 587972 218540 595672 218568
rect 587972 218484 588028 218540
rect 459442 218428 459452 218484
rect 459508 218428 588028 218484
rect -960 206164 480 206360
rect -960 206136 532 206164
rect 392 206108 532 206136
rect 476 206052 532 206108
rect 364 205996 532 206052
rect 364 205044 420 205996
rect 595560 205380 597000 205576
rect 587972 205352 597000 205380
rect 587972 205324 595672 205352
rect 587972 205044 588028 205324
rect 364 204988 52892 205044
rect 52948 204988 52958 205044
rect 446002 204988 446012 205044
rect 446068 204988 588028 205044
rect 590482 192332 590492 192388
rect 590548 192360 595672 192388
rect 590548 192332 597000 192360
rect -960 192052 480 192248
rect 595560 192136 597000 192332
rect -960 192024 532 192052
rect 392 191996 532 192024
rect 476 191940 532 191996
rect 364 191884 532 191940
rect 364 191604 420 191884
rect 364 191548 22652 191604
rect 22708 191548 22718 191604
rect 595560 178948 597000 179144
rect 595420 178920 597000 178948
rect 595420 178892 595672 178920
rect 595420 178836 595476 178892
rect 595420 178780 595700 178836
rect 595644 178164 595700 178780
rect -960 177940 480 178136
rect 454402 178108 454412 178164
rect 454468 178108 595700 178164
rect -960 177912 532 177940
rect 392 177884 532 177912
rect 476 177828 532 177884
rect 364 177772 532 177828
rect 364 176484 420 177772
rect 364 176428 29372 176484
rect 29428 176428 29438 176484
rect 593842 165900 593852 165956
rect 593908 165928 595672 165956
rect 593908 165900 597000 165928
rect 595560 165704 597000 165900
rect -960 163828 480 164024
rect -960 163800 532 163828
rect 392 163772 532 163800
rect 476 163716 532 163772
rect 364 163660 532 163716
rect 364 163044 420 163660
rect 364 162988 51212 163044
rect 51268 162988 51278 163044
rect 593730 152684 593740 152740
rect 593796 152712 595672 152740
rect 593796 152684 597000 152712
rect 595560 152488 597000 152684
rect -960 149716 480 149912
rect -960 149688 11788 149716
rect 392 149660 11788 149688
rect 11732 149604 11788 149660
rect 11732 149548 27692 149604
rect 27748 149548 27758 149604
rect 595560 139300 597000 139496
rect 595420 139272 597000 139300
rect 595420 139244 595672 139272
rect 595420 139188 595476 139244
rect 595420 139132 595700 139188
rect 595644 137844 595700 139132
rect 477922 137788 477932 137844
rect 477988 137788 595700 137844
rect -960 135604 480 135800
rect -960 135576 532 135604
rect 392 135548 532 135576
rect 476 135492 532 135548
rect 364 135436 532 135492
rect 364 134484 420 135436
rect 364 134428 32732 134484
rect 32788 134428 32798 134484
rect 593618 126252 593628 126308
rect 593684 126280 595672 126308
rect 593684 126252 597000 126280
rect 595560 126056 597000 126252
rect 392 121688 9212 121716
rect -960 121660 9212 121688
rect 9268 121660 9278 121716
rect -960 121464 480 121660
rect 595560 112868 597000 113064
rect 587972 112840 597000 112868
rect 587972 112812 595672 112840
rect 587972 112644 588028 112812
rect 456082 112588 456092 112644
rect 456148 112588 588028 112644
rect -960 107492 480 107576
rect -960 107436 2492 107492
rect 2548 107436 2558 107492
rect -960 107352 480 107436
rect 595560 99652 597000 99848
rect 595420 99624 597000 99652
rect 595420 99596 595672 99624
rect 595420 99540 595476 99596
rect 595420 99484 595700 99540
rect 595644 99204 595700 99484
rect 476242 99148 476252 99204
rect 476308 99148 595700 99204
rect -960 93268 480 93464
rect -960 93240 532 93268
rect 392 93212 532 93240
rect 476 93156 532 93212
rect 364 93100 532 93156
rect 364 92484 420 93100
rect 364 92428 17612 92484
rect 17668 92428 17678 92484
rect 593506 86604 593516 86660
rect 593572 86632 595672 86660
rect 593572 86604 597000 86632
rect 595560 86408 597000 86604
rect -960 79156 480 79352
rect -960 79128 11788 79156
rect 392 79100 11788 79128
rect 11732 79044 11788 79100
rect 11732 78988 49532 79044
rect 49588 78988 49598 79044
rect 593394 73388 593404 73444
rect 593460 73416 595672 73444
rect 593460 73388 597000 73416
rect 595560 73192 597000 73388
rect -960 65044 480 65240
rect -960 65016 532 65044
rect 392 64988 532 65016
rect 476 64932 532 64988
rect 364 64876 532 64932
rect 364 63924 420 64876
rect 364 63868 44492 63924
rect 44548 63868 44558 63924
rect 595560 60004 597000 60200
rect 595420 59976 597000 60004
rect 595420 59948 595672 59976
rect 595420 59892 595476 59948
rect 595420 59836 595700 59892
rect 90738 59388 90748 59444
rect 90804 59388 91644 59444
rect 91700 59388 91710 59444
rect 109218 59388 109228 59444
rect 109284 59388 110124 59444
rect 110180 59388 110190 59444
rect 114258 59388 114268 59444
rect 114324 59388 115052 59444
rect 115108 59388 115118 59444
rect 142818 59388 142828 59444
rect 142884 59388 143388 59444
rect 143444 59388 143454 59444
rect 146178 59388 146188 59444
rect 146244 59388 147084 59444
rect 147140 59388 147150 59444
rect 193218 59388 193228 59444
rect 193284 59388 193900 59444
rect 193956 59388 193966 59444
rect 220098 59388 220108 59444
rect 220164 59388 221004 59444
rect 221060 59388 221070 59444
rect 238578 59388 238588 59444
rect 238644 59388 239484 59444
rect 239540 59388 239550 59444
rect 294018 59388 294028 59444
rect 294084 59388 294924 59444
rect 294980 59388 294990 59444
rect 312498 59388 312508 59444
rect 312564 59388 313404 59444
rect 313460 59388 313470 59444
rect 341058 59388 341068 59444
rect 341124 59388 341740 59444
rect 341796 59388 341806 59444
rect 349458 59388 349468 59444
rect 349524 59388 350364 59444
rect 350420 59388 350430 59444
rect 386418 59388 386428 59444
rect 386484 59388 387324 59444
rect 387380 59388 387390 59444
rect 433458 59388 433468 59444
rect 433524 59388 434140 59444
rect 434196 59388 434206 59444
rect 290658 59276 290668 59332
rect 290724 59276 291228 59332
rect 291284 59276 291294 59332
rect 304098 59052 304108 59108
rect 304164 59052 304780 59108
rect 304836 59052 304846 59108
rect 595644 58884 595700 59836
rect 496402 58828 496412 58884
rect 496468 58828 595700 58884
rect 354610 58044 354620 58100
rect 354676 58044 458668 58100
rect 458724 58044 458734 58100
rect 378130 57932 378140 57988
rect 378196 57932 493948 57988
rect 494004 57932 494024 57988
rect 258738 56812 258748 56868
rect 258804 56812 264572 56868
rect 264628 56812 264638 56868
rect 344418 56812 344428 56868
rect 344484 56812 355292 56868
rect 355348 56812 355358 56868
rect 366258 56812 366268 56868
rect 366324 56812 372092 56868
rect 372148 56812 372158 56868
rect 426738 56812 426748 56868
rect 426804 56812 446012 56868
rect 446068 56812 446078 56868
rect 91522 56700 91532 56756
rect 91588 56700 95788 56756
rect 95844 56700 95854 56756
rect 98690 56700 98700 56756
rect 98756 56700 107548 56756
rect 107604 56700 107614 56756
rect 236898 56700 236908 56756
rect 236964 56700 242732 56756
rect 242788 56700 242798 56756
rect 255378 56700 255388 56756
rect 255444 56700 261212 56756
rect 261268 56700 261278 56756
rect 285730 56700 285740 56756
rect 285796 56700 325052 56756
rect 325108 56700 325118 56756
rect 325938 56700 325948 56756
rect 326004 56700 330092 56756
rect 330148 56700 330158 56756
rect 331202 56700 331212 56756
rect 331268 56700 351932 56756
rect 351988 56700 351998 56756
rect 384738 56700 384748 56756
rect 384804 56700 390348 56756
rect 390404 56700 390414 56756
rect 393138 56700 393148 56756
rect 393204 56700 412412 56756
rect 412468 56700 412478 56756
rect 431778 56700 431788 56756
rect 431844 56700 454412 56756
rect 454468 56700 454478 56756
rect 62962 56588 62972 56644
rect 63028 56588 72268 56644
rect 72324 56588 72334 56644
rect 83122 56588 83132 56644
rect 83188 56588 100828 56644
rect 100884 56588 100894 56644
rect 140242 56588 140252 56644
rect 140308 56588 146188 56644
rect 146244 56588 146254 56644
rect 221778 56588 221788 56644
rect 221844 56588 227612 56644
rect 227668 56588 227678 56644
rect 290882 56588 290892 56644
rect 290948 56588 296492 56644
rect 296548 56588 296558 56644
rect 317650 56588 317660 56644
rect 317716 56588 370412 56644
rect 370468 56588 370478 56644
rect 383170 56588 383180 56644
rect 383236 56588 393596 56644
rect 393652 56588 393662 56644
rect 398178 56588 398188 56644
rect 398244 56588 444332 56644
rect 444388 56588 444398 56644
rect 68002 56476 68012 56532
rect 68068 56476 95900 56532
rect 95956 56476 95966 56532
rect 99922 56476 99932 56532
rect 99988 56476 109228 56532
rect 109284 56476 109294 56532
rect 135202 56476 135212 56532
rect 135268 56476 142828 56532
rect 142884 56476 142894 56532
rect 203298 56476 203308 56532
rect 203364 56476 210812 56532
rect 210868 56476 210878 56532
rect 211810 56476 211820 56532
rect 211876 56476 229292 56532
rect 229348 56476 229358 56532
rect 248770 56476 248780 56532
rect 248836 56476 266252 56532
rect 266308 56476 266318 56532
rect 267250 56476 267260 56532
rect 267316 56476 279692 56532
rect 279748 56476 279758 56532
rect 290658 56476 290668 56532
rect 290724 56476 356972 56532
rect 357028 56476 357038 56532
rect 364690 56476 364700 56532
rect 364756 56476 432572 56532
rect 432628 56476 432638 56532
rect 56242 56364 56252 56420
rect 56308 56364 90748 56420
rect 90804 56364 90814 56420
rect 107538 56364 107548 56420
rect 107604 56364 127708 56420
rect 127764 56364 127774 56420
rect 128482 56364 128492 56420
rect 128548 56364 132748 56420
rect 132804 56364 132814 56420
rect 136210 56364 136220 56420
rect 136276 56364 146300 56420
rect 146356 56364 146366 56420
rect 171602 56364 171612 56420
rect 171668 56364 176428 56420
rect 176484 56364 176494 56420
rect 210018 56364 210028 56420
rect 210084 56364 214172 56420
rect 214228 56364 214238 56420
rect 218418 56364 218428 56420
rect 218484 56364 224252 56420
rect 224308 56364 224318 56420
rect 225250 56364 225260 56420
rect 225316 56364 251132 56420
rect 251188 56364 251198 56420
rect 253810 56364 253820 56420
rect 253876 56364 286412 56420
rect 286468 56364 286478 56420
rect 294018 56364 294028 56420
rect 294084 56364 362012 56420
rect 362068 56364 362078 56420
rect 362898 56364 362908 56420
rect 362964 56364 365596 56420
rect 365652 56364 365662 56420
rect 386530 56364 386540 56420
rect 386596 56364 484652 56420
rect 484708 56364 484718 56420
rect 28578 56252 28588 56308
rect 28644 56252 75628 56308
rect 75684 56252 75694 56308
rect 94882 56252 94892 56308
rect 94948 56252 115948 56308
rect 116004 56252 116014 56308
rect 125122 56252 125132 56308
rect 125188 56252 137788 56308
rect 137844 56252 137854 56308
rect 174850 56252 174860 56308
rect 174916 56252 180572 56308
rect 180628 56252 180638 56308
rect 184818 56252 184828 56308
rect 184884 56252 190652 56308
rect 190708 56252 190718 56308
rect 213378 56252 213388 56308
rect 213444 56252 234332 56308
rect 234388 56252 234398 56308
rect 235330 56252 235340 56308
rect 235396 56252 267932 56308
rect 267988 56252 267998 56308
rect 275650 56252 275660 56308
rect 275716 56252 335132 56308
rect 335188 56252 335198 56308
rect 336130 56252 336140 56308
rect 336196 56252 427532 56308
rect 427588 56252 427598 56308
rect 428418 56252 428428 56308
rect 428484 56252 570332 56308
rect 570388 56252 570398 56308
rect 309362 55804 309372 55860
rect 309428 55804 315980 55860
rect 316036 55804 316046 55860
rect 144498 55580 144508 55636
rect 144564 55580 151340 55636
rect 151396 55580 151406 55636
rect 199938 55580 199948 55636
rect 200004 55580 202412 55636
rect 202468 55580 202478 55636
rect 76402 55468 76412 55524
rect 76468 55468 77308 55524
rect 77364 55468 77374 55524
rect 84802 55468 84812 55524
rect 84868 55468 87388 55524
rect 87444 55468 87454 55524
rect 89170 55468 89180 55524
rect 89236 55468 92428 55524
rect 92484 55468 92494 55524
rect 110002 55468 110012 55524
rect 110068 55468 110908 55524
rect 110964 55468 110974 55524
rect 113362 55468 113372 55524
rect 113428 55468 114268 55524
rect 114324 55468 114334 55524
rect 114482 55468 114492 55524
rect 114548 55468 116060 55524
rect 116116 55468 116126 55524
rect 118402 55468 118412 55524
rect 118468 55468 119308 55524
rect 119364 55468 119374 55524
rect 123442 55468 123452 55524
rect 123508 55468 124348 55524
rect 124404 55468 124414 55524
rect 131842 55468 131852 55524
rect 131908 55468 134428 55524
rect 134484 55468 134494 55524
rect 135426 55468 135436 55524
rect 135492 55468 136108 55524
rect 136164 55468 136174 55524
rect 148642 55468 148652 55524
rect 148708 55468 151228 55524
rect 151284 55468 151294 55524
rect 164770 55468 164780 55524
rect 164836 55468 166460 55524
rect 166516 55468 166526 55524
rect 168018 55468 168028 55524
rect 168084 55468 171388 55524
rect 171444 55468 171454 55524
rect 176642 55468 176652 55524
rect 176708 55468 178892 55524
rect 178948 55468 178958 55524
rect 183250 55468 183260 55524
rect 183316 55468 185612 55524
rect 185668 55468 185678 55524
rect 201730 55468 201740 55524
rect 201796 55468 204092 55524
rect 204148 55468 204158 55524
rect 206770 55468 206780 55524
rect 206836 55468 209132 55524
rect 209188 55468 209198 55524
rect 240258 55468 240268 55524
rect 240324 55468 246092 55524
rect 246148 55468 246158 55524
rect 272290 55468 272300 55524
rect 272356 55468 274652 55524
rect 274708 55468 274718 55524
rect 294242 55468 294252 55524
rect 294308 55468 298172 55524
rect 298228 55468 298238 55524
rect 309138 55468 309148 55524
rect 309204 55468 311612 55524
rect 311668 55468 311678 55524
rect 312610 55468 312620 55524
rect 312676 55468 314972 55524
rect 315028 55468 315038 55524
rect 330978 55468 330988 55524
rect 331044 55468 333452 55524
rect 333508 55468 333518 55524
rect 381378 55468 381388 55524
rect 381444 55468 383852 55524
rect 383908 55468 383918 55524
rect 391570 55468 391580 55524
rect 391636 55468 393932 55524
rect 393988 55468 393998 55524
rect 401650 55468 401660 55524
rect 401716 55468 407372 55524
rect 407428 55468 407438 55524
rect 347778 54908 347788 54964
rect 347844 54908 448588 54964
rect 448644 54908 448654 54964
rect 53778 54796 53788 54852
rect 53844 54796 89180 54852
rect 89236 54796 89246 54852
rect 410050 54796 410060 54852
rect 410116 54796 544348 54852
rect 544404 54796 544414 54852
rect 36082 54684 36092 54740
rect 36148 54684 78988 54740
rect 79044 54684 79054 54740
rect 278898 54684 278908 54740
rect 278964 54684 342748 54740
rect 342804 54684 342814 54740
rect 416658 54684 416668 54740
rect 416724 54684 554428 54740
rect 554484 54684 554494 54740
rect 36978 54572 36988 54628
rect 37044 54572 82460 54628
rect 82516 54572 82526 54628
rect 312498 54572 312508 54628
rect 312564 54572 394828 54628
rect 394884 54572 394894 54628
rect 420130 54572 420140 54628
rect 420196 54572 560252 54628
rect 560308 54572 560318 54628
rect 77298 53116 77308 53172
rect 77364 53116 98700 53172
rect 98756 53116 98766 53172
rect 349570 53116 349580 53172
rect 349636 53116 450268 53172
rect 450324 53116 450334 53172
rect 34514 53004 34524 53060
rect 34580 53004 73948 53060
rect 74004 53004 74014 53060
rect 373090 53004 373100 53060
rect 373156 53004 487228 53060
rect 487284 53004 487294 53060
rect 31938 52892 31948 52948
rect 32004 52892 77420 52948
rect 77476 52892 77486 52948
rect 423490 52892 423500 52948
rect 423556 52892 566188 52948
rect 566244 52892 566254 52948
rect 359650 51436 359660 51492
rect 359716 51436 465388 51492
rect 465444 51436 465454 51492
rect 365586 51324 365596 51380
rect 365652 51324 472108 51380
rect 472164 51324 472174 51380
rect 40338 51212 40348 51268
rect 40404 51212 84028 51268
rect 84084 51212 84094 51268
rect 396610 51212 396620 51268
rect 396676 51212 522508 51268
rect 522564 51212 522574 51268
rect -960 50932 480 51128
rect -960 50904 532 50932
rect 392 50876 532 50904
rect 476 50820 532 50876
rect 364 50764 532 50820
rect 364 50484 420 50764
rect 364 50428 34412 50484
rect 34468 50428 34478 50484
rect 390338 49644 390348 49700
rect 390404 49644 505708 49700
rect 505764 49644 505774 49700
rect 315970 49532 315980 49588
rect 316036 49532 389788 49588
rect 389844 49532 389854 49588
rect 403218 49532 403228 49588
rect 403284 49532 534268 49588
rect 534324 49532 534334 49588
rect 356178 48076 356188 48132
rect 356244 48076 462028 48132
rect 462084 48076 462094 48132
rect 310818 47964 310828 48020
rect 310884 47964 391580 48020
rect 391636 47964 391646 48020
rect 393586 47964 393596 48020
rect 393652 47964 502348 48020
rect 502404 47964 502414 48020
rect 238690 47852 238700 47908
rect 238756 47852 278908 47908
rect 278964 47852 278974 47908
rect 389890 47852 389900 47908
rect 389956 47852 514108 47908
rect 514164 47852 514174 47908
rect 593282 46956 593292 47012
rect 593348 46984 595672 47012
rect 593348 46956 597000 46984
rect 595560 46760 597000 46956
rect 342850 46396 342860 46452
rect 342916 46396 440300 46452
rect 440356 46396 440366 46452
rect 368050 46284 368060 46340
rect 368116 46284 480508 46340
rect 480564 46284 480574 46340
rect 299170 46172 299180 46228
rect 299236 46172 374780 46228
rect 374836 46172 374846 46228
rect 383842 46172 383852 46228
rect 383908 46172 500668 46228
rect 500724 46172 500734 46228
rect 346210 44716 346220 44772
rect 346276 44716 446908 44772
rect 446964 44716 446984 44772
rect 393922 44604 393932 44660
rect 393988 44604 515788 44660
rect 515844 44604 515854 44660
rect 58818 44492 58828 44548
rect 58884 44492 91532 44548
rect 91588 44492 91598 44548
rect 265458 44492 265468 44548
rect 265524 44492 320908 44548
rect 320964 44492 320974 44548
rect 321122 44492 321132 44548
rect 321188 44492 406588 44548
rect 406644 44492 406654 44548
rect 407362 44492 407372 44548
rect 407428 44492 530908 44548
rect 530964 44492 530974 44548
rect 372082 42924 372092 42980
rect 372148 42924 477148 42980
rect 477204 42924 477214 42980
rect 60386 42812 60396 42868
rect 60452 42812 590492 42868
rect 590548 42812 590558 42868
rect 357858 41356 357868 41412
rect 357924 41356 463708 41412
rect 463764 41356 463774 41412
rect 415090 41244 415100 41300
rect 415156 41244 551068 41300
rect 551124 41244 551134 41300
rect 4946 41132 4956 41188
rect 5012 41132 440188 41188
rect 440244 41132 440254 41188
rect 359538 39564 359548 39620
rect 359604 39564 467068 39620
rect 467124 39564 467134 39620
rect 334338 39452 334348 39508
rect 334404 39452 428428 39508
rect 428484 39452 428494 39508
rect 446002 39452 446012 39508
rect 446068 39452 571228 39508
rect 571284 39452 571294 39508
rect 333442 37996 333452 38052
rect 333508 37996 421708 38052
rect 421764 37996 421774 38052
rect 388322 37884 388332 37940
rect 388388 37884 512428 37940
rect 512484 37884 512494 37940
rect 264562 37772 264572 37828
rect 264628 37772 310828 37828
rect 310884 37772 310894 37828
rect 311602 37772 311612 37828
rect 311668 37772 388108 37828
rect 388164 37772 388174 37828
rect 401538 37772 401548 37828
rect 401604 37772 532588 37828
rect 532644 37772 532654 37828
rect -960 36932 480 37016
rect -960 36876 4956 36932
rect 5012 36876 5022 36932
rect -960 36792 480 36876
rect 19282 36204 19292 36260
rect 19348 36204 69020 36260
rect 69076 36204 69086 36260
rect 354498 36204 354508 36260
rect 354564 36204 460348 36260
rect 460404 36204 460414 36260
rect 15138 36092 15148 36148
rect 15204 36092 67228 36148
rect 67284 36092 67294 36148
rect 243730 36092 243740 36148
rect 243796 36092 288988 36148
rect 289044 36092 289054 36148
rect 314962 36092 314972 36148
rect 315028 36092 393148 36148
rect 393204 36092 393214 36148
rect 421810 36092 421820 36148
rect 421876 36092 562828 36148
rect 562884 36092 562894 36148
rect 346098 34524 346108 34580
rect 346164 34524 445228 34580
rect 445284 34524 445294 34580
rect 261202 34412 261212 34468
rect 261268 34412 305900 34468
rect 305956 34412 305966 34468
rect 374658 34412 374668 34468
rect 374724 34412 490588 34468
rect 490644 34412 490654 34468
rect 593170 33740 593180 33796
rect 593236 33768 595672 33796
rect 593236 33740 597000 33768
rect 595560 33544 597000 33740
rect 327730 32844 327740 32900
rect 327796 32844 418460 32900
rect 418516 32844 418526 32900
rect 454402 32844 454412 32900
rect 454468 32844 579628 32900
rect 579684 32844 579694 32900
rect 274642 32732 274652 32788
rect 274708 32732 332780 32788
rect 332836 32732 332846 32788
rect 394930 32732 394940 32788
rect 394996 32732 520828 32788
rect 520884 32732 520894 32788
rect 298162 31164 298172 31220
rect 298228 31164 364700 31220
rect 364756 31164 364766 31220
rect 371298 31164 371308 31220
rect 371364 31164 485548 31220
rect 485604 31164 485614 31220
rect 322690 31052 322700 31108
rect 322756 31052 408380 31108
rect 408436 31052 408446 31108
rect 428530 31052 428540 31108
rect 428596 31052 574588 31108
rect 574644 31052 574654 31108
rect 277218 29484 277228 29540
rect 277284 29484 339500 29540
rect 339556 29484 339566 29540
rect 351138 29484 351148 29540
rect 351204 29484 453628 29540
rect 453684 29484 453694 29540
rect 224242 29372 224252 29428
rect 224308 29372 248780 29428
rect 248836 29372 248846 29428
rect 280690 29372 280700 29428
rect 280756 29372 346108 29428
rect 346164 29372 346174 29428
rect 369618 29372 369628 29428
rect 369684 29372 482188 29428
rect 482244 29372 482254 29428
rect 296482 27804 296492 27860
rect 296548 27804 359548 27860
rect 359604 27804 359614 27860
rect 406690 27804 406700 27860
rect 406756 27804 539308 27860
rect 539364 27804 539374 27860
rect 44482 27692 44492 27748
rect 44548 27692 82348 27748
rect 82404 27692 82414 27748
rect 317538 27692 317548 27748
rect 317604 27692 403228 27748
rect 403284 27692 403294 27748
rect 425058 27692 425068 27748
rect 425124 27692 567868 27748
rect 567924 27692 567934 27748
rect 289090 26124 289100 26180
rect 289156 26124 357868 26180
rect 357924 26124 357934 26180
rect 367938 26124 367948 26180
rect 368004 26124 478828 26180
rect 478884 26124 478894 26180
rect 48738 26012 48748 26068
rect 48804 26012 89068 26068
rect 89124 26012 89134 26068
rect 230290 26012 230300 26068
rect 230356 26012 265468 26068
rect 265524 26012 265534 26068
rect 304210 26012 304220 26068
rect 304276 26012 379820 26068
rect 379876 26012 379886 26068
rect 418338 26012 418348 26068
rect 418404 26012 557788 26068
rect 557844 26012 557854 26068
rect 52098 25116 52108 25172
rect 52164 25116 56252 25172
rect 56308 25116 56318 25172
rect 307458 24556 307468 24612
rect 307524 24556 386540 24612
rect 386596 24556 386606 24612
rect 383058 24444 383068 24500
rect 383124 24444 504028 24500
rect 504084 24444 504094 24500
rect 257170 24332 257180 24388
rect 257236 24332 308252 24388
rect 308308 24332 308318 24388
rect 386418 24332 386428 24388
rect 386484 24332 509068 24388
rect 509124 24332 509134 24388
rect -960 22708 480 22904
rect 332658 22764 332668 22820
rect 332724 22764 425068 22820
rect 425124 22764 425134 22820
rect -960 22680 532 22708
rect 392 22652 532 22680
rect 10098 22652 10108 22708
rect 10164 22652 63868 22708
rect 63924 22652 63934 22708
rect 379698 22652 379708 22708
rect 379764 22652 497308 22708
rect 497364 22652 497374 22708
rect 476 22596 532 22652
rect 364 22540 532 22596
rect 364 21924 420 22540
rect 364 21868 436828 21924
rect 436884 21868 436894 21924
rect 341170 21084 341180 21140
rect 341236 21084 436828 21140
rect 436884 21084 436894 21140
rect 30258 20972 30268 21028
rect 30324 20972 76412 21028
rect 76468 20972 76478 21028
rect 82338 20972 82348 21028
rect 82404 20972 110012 21028
rect 110068 20972 110078 21028
rect 246082 20972 246092 21028
rect 246148 20972 282380 21028
rect 282436 20972 282446 21028
rect 361218 20972 361228 21028
rect 361284 20972 468748 21028
rect 468804 20972 468814 21028
rect 590482 20524 590492 20580
rect 590548 20552 595672 20580
rect 590548 20524 597000 20552
rect 595560 20328 597000 20524
rect 297378 19516 297388 19572
rect 297444 19516 371308 19572
rect 371364 19516 371374 19572
rect 352818 19404 352828 19460
rect 352884 19404 456092 19460
rect 456148 19404 456158 19460
rect 47058 19292 47068 19348
rect 47124 19292 87500 19348
rect 87556 19292 87566 19348
rect 250338 19292 250348 19348
rect 250404 19292 297388 19348
rect 297444 19292 297454 19348
rect 314178 19292 314188 19348
rect 314244 19292 396620 19348
rect 396676 19292 396686 19348
rect 405010 19292 405020 19348
rect 405076 19292 537628 19348
rect 537684 19292 537694 19348
rect 241938 17948 241948 18004
rect 242004 17948 285740 18004
rect 285796 17948 285806 18004
rect 325042 17948 325052 18004
rect 325108 17948 352828 18004
rect 352884 17948 352904 18004
rect 351922 17836 351932 17892
rect 351988 17836 423500 17892
rect 423556 17836 423566 17892
rect 432562 17836 432572 17892
rect 432628 17836 475468 17892
rect 475524 17836 475534 17892
rect 285618 17724 285628 17780
rect 285684 17724 351148 17780
rect 351204 17724 351214 17780
rect 355282 17724 355292 17780
rect 355348 17724 443548 17780
rect 443604 17724 443614 17780
rect 45378 17612 45388 17668
rect 45444 17612 84812 17668
rect 84868 17612 84878 17668
rect 242722 17612 242732 17668
rect 242788 17612 277228 17668
rect 277284 17612 277294 17668
rect 295698 17612 295708 17668
rect 295764 17612 367948 17668
rect 368004 17612 368014 17668
rect 396498 17612 396508 17668
rect 396564 17612 523292 17668
rect 523348 17612 523358 17668
rect 209122 16156 209132 16212
rect 209188 16156 231980 16212
rect 232036 16156 232046 16212
rect 75618 16044 75628 16100
rect 75684 16044 105980 16100
rect 106036 16044 106046 16100
rect 220210 16044 220220 16100
rect 220276 16044 250348 16100
rect 250404 16044 250414 16100
rect 267138 16044 267148 16100
rect 267204 16044 322700 16100
rect 322756 16044 322766 16100
rect 349458 16044 349468 16100
rect 349524 16044 451948 16100
rect 452004 16044 452014 16100
rect 63858 15932 63868 15988
rect 63924 15932 99148 15988
rect 99204 15932 99214 15988
rect 115938 15932 115948 15988
rect 116004 15932 128492 15988
rect 128548 15932 128558 15988
rect 231858 15932 231868 15988
rect 231924 15932 268940 15988
rect 268996 15932 269006 15988
rect 305778 15932 305788 15988
rect 305844 15932 383068 15988
rect 383124 15932 383134 15988
rect 413298 15932 413308 15988
rect 413364 15932 549388 15988
rect 549444 15932 549454 15988
rect 220098 14588 220108 14644
rect 220164 14588 252140 14644
rect 252196 14588 252206 14644
rect 315858 14588 315868 14644
rect 315924 14588 399980 14644
rect 400036 14588 400046 14644
rect 252018 14364 252028 14420
rect 252084 14364 300860 14420
rect 300916 14364 300926 14420
rect 399858 14364 399868 14420
rect 399924 14364 529228 14420
rect 529284 14364 529294 14420
rect 69010 14252 69020 14308
rect 69076 14252 102508 14308
rect 102564 14252 102574 14308
rect 102722 14252 102732 14308
rect 102788 14252 124460 14308
rect 124516 14252 124526 14308
rect 202402 14252 202412 14308
rect 202468 14252 220108 14308
rect 220164 14252 220174 14308
rect 262210 14252 262220 14308
rect 262276 14252 315868 14308
rect 315924 14252 315934 14308
rect 322578 14252 322588 14308
rect 322644 14252 410060 14308
rect 410116 14252 410126 14308
rect 433570 14252 433580 14308
rect 433636 14252 581308 14308
rect 581364 14252 581374 14308
rect 273858 12796 273868 12852
rect 273924 12796 334348 12852
rect 334404 12796 334414 12852
rect 337698 12796 337708 12852
rect 337764 12796 433580 12852
rect 433636 12796 433646 12852
rect 27682 12684 27692 12740
rect 27748 12684 72716 12740
rect 72772 12684 72782 12740
rect 198370 12684 198380 12740
rect 198436 12684 215852 12740
rect 215908 12684 215918 12740
rect 238578 12684 238588 12740
rect 238644 12684 280700 12740
rect 280756 12684 280766 12740
rect 299058 12684 299068 12740
rect 299124 12684 374668 12740
rect 374724 12684 374734 12740
rect 414978 12684 414988 12740
rect 415044 12684 552748 12740
rect 552804 12684 552814 12740
rect 72482 12572 72492 12628
rect 72548 12572 104188 12628
rect 104244 12572 104254 12628
rect 104402 12572 104412 12628
rect 104468 12572 123452 12628
rect 123508 12572 123518 12628
rect 215058 12572 215068 12628
rect 215124 12572 243740 12628
rect 243796 12572 243806 12628
rect 268818 12572 268828 12628
rect 268884 12572 325948 12628
rect 326004 12572 326014 12628
rect 327618 12572 327628 12628
rect 327684 12572 415772 12628
rect 415828 12572 415838 12628
rect 430098 12572 430108 12628
rect 430164 12572 576268 12628
rect 576324 12572 576334 12628
rect 216850 11340 216860 11396
rect 216916 11340 247436 11396
rect 247492 11340 247502 11396
rect 246978 11116 246988 11172
rect 247044 11116 293132 11172
rect 293188 11116 293198 11172
rect 319218 11116 319228 11172
rect 319284 11116 405468 11172
rect 405524 11116 405534 11172
rect 270498 11004 270508 11060
rect 270564 11004 329308 11060
rect 329364 11004 329384 11060
rect 336018 11004 336028 11060
rect 336084 11004 432124 11060
rect 432180 11004 432190 11060
rect 22978 10892 22988 10948
rect 23044 10892 62972 10948
rect 63028 10892 63038 10948
rect 89618 10892 89628 10948
rect 89684 10892 113372 10948
rect 113428 10892 113438 10948
rect 198258 10892 198268 10948
rect 198324 10892 218316 10948
rect 218372 10892 218382 10948
rect 225138 10892 225148 10948
rect 225204 10892 260764 10948
rect 260820 10892 260830 10948
rect 287298 10892 287308 10948
rect 287364 10892 355964 10948
rect 356020 10892 356030 10948
rect 391458 10892 391468 10948
rect 391524 10892 517804 10948
rect 517860 10892 517870 10948
rect 570322 10108 570332 10164
rect 570388 10108 573020 10164
rect 573076 10108 573086 10164
rect 216738 9324 216748 9380
rect 216804 9324 245532 9380
rect 245588 9324 245598 9380
rect 330082 9324 330092 9380
rect 330148 9324 414988 9380
rect 415044 9324 415054 9380
rect 444322 9324 444332 9380
rect 444388 9324 527324 9380
rect 527380 9324 527390 9380
rect 120082 9212 120092 9268
rect 120148 9212 131852 9268
rect 131908 9212 131918 9268
rect 235218 9212 235228 9268
rect 235284 9212 274092 9268
rect 274148 9212 274158 9268
rect 279682 9212 279692 9268
rect 279748 9212 325500 9268
rect 325556 9212 325566 9268
rect 378018 9212 378028 9268
rect 378084 9212 496860 9268
rect 496916 9212 496926 9268
rect -960 8596 480 8792
rect -960 8568 11788 8596
rect 392 8540 11788 8568
rect 11732 8484 11788 8540
rect 11732 8428 441868 8484
rect 441924 8428 441934 8484
rect 356962 8092 356972 8148
rect 357028 8092 361676 8148
rect 361732 8092 361742 8148
rect 142706 7980 142716 8036
rect 142772 7980 144732 8036
rect 144788 7980 144798 8036
rect 286402 7868 286412 7924
rect 286468 7868 304556 7924
rect 304612 7868 304622 7924
rect 370402 7868 370412 7924
rect 370468 7868 401660 7924
rect 401716 7868 401726 7924
rect 82002 7756 82012 7812
rect 82068 7756 99932 7812
rect 99988 7756 99998 7812
rect 196578 7756 196588 7812
rect 196644 7756 215068 7812
rect 215124 7756 215134 7812
rect 266242 7756 266252 7812
rect 266308 7756 296940 7812
rect 296996 7756 297006 7812
rect 302418 7756 302428 7812
rect 302484 7756 378812 7812
rect 378868 7756 378878 7812
rect 411572 7756 413084 7812
rect 413140 7756 413150 7812
rect 411572 7700 411628 7756
rect 99026 7644 99036 7700
rect 99092 7644 120988 7700
rect 121044 7644 121054 7700
rect 132626 7644 132636 7700
rect 132692 7644 141148 7700
rect 141204 7644 141224 7700
rect 214162 7644 214172 7700
rect 214228 7644 236012 7700
rect 236068 7644 236078 7700
rect 243618 7644 243628 7700
rect 243684 7644 287420 7700
rect 287476 7644 287486 7700
rect 324258 7644 324268 7700
rect 324324 7644 411628 7700
rect 412402 7644 412412 7700
rect 412468 7644 519708 7700
rect 519764 7644 519774 7700
rect 36306 7532 36316 7588
rect 36372 7532 80668 7588
rect 80724 7532 80734 7588
rect 95330 7532 95340 7588
rect 95396 7532 118412 7588
rect 118468 7532 118478 7588
rect 121986 7532 121996 7588
rect 122052 7532 135436 7588
rect 135492 7532 135502 7588
rect 137778 7532 137788 7588
rect 137844 7532 143276 7588
rect 143332 7532 143342 7588
rect 152450 7532 152460 7588
rect 152516 7532 156380 7588
rect 156436 7532 156446 7588
rect 181458 7532 181468 7588
rect 181524 7532 192220 7588
rect 192276 7532 192286 7588
rect 204082 7532 204092 7588
rect 204148 7532 224588 7588
rect 224644 7532 224654 7588
rect 228498 7532 228508 7588
rect 228564 7532 264572 7588
rect 264628 7532 264638 7588
rect 283938 7532 283948 7588
rect 284004 7532 350252 7588
rect 350308 7532 350318 7588
rect 372978 7532 372988 7588
rect 373044 7532 489244 7588
rect 489300 7532 489310 7588
rect 594290 7308 594300 7364
rect 594356 7336 595672 7364
rect 594356 7308 597000 7336
rect 595560 7112 597000 7308
rect 142930 6748 142940 6804
rect 142996 6748 149548 6804
rect 149604 6748 149614 6804
rect 427522 6748 427532 6804
rect 427588 6748 430220 6804
rect 430276 6748 430286 6804
rect 190642 6300 190652 6356
rect 190708 6300 197932 6356
rect 197988 6300 197998 6356
rect 362002 6300 362012 6356
rect 362068 6300 367388 6356
rect 367444 6300 367454 6356
rect 185602 6188 185612 6244
rect 185668 6188 196028 6244
rect 196084 6188 196094 6244
rect 234322 6188 234332 6244
rect 234388 6188 241724 6244
rect 241780 6188 241790 6244
rect 260418 6188 260428 6244
rect 260484 6188 314188 6244
rect 314244 6188 314254 6244
rect 329410 6188 329420 6244
rect 329476 6188 420700 6244
rect 420756 6188 420766 6244
rect 91522 6076 91532 6132
rect 91588 6076 94892 6132
rect 94948 6076 94958 6132
rect 110562 6076 110572 6132
rect 110628 6076 127820 6132
rect 127876 6076 127886 6132
rect 210802 6076 210812 6132
rect 210868 6076 226492 6132
rect 226548 6076 226558 6132
rect 229282 6076 229292 6132
rect 229348 6076 237916 6132
rect 237972 6076 237982 6132
rect 251122 6076 251132 6132
rect 251188 6076 258860 6132
rect 258916 6076 258926 6132
rect 262098 6076 262108 6132
rect 262164 6076 317884 6132
rect 317940 6076 317950 6132
rect 341058 6076 341068 6132
rect 341124 6076 439740 6132
rect 439796 6076 439806 6132
rect 61058 5964 61068 6020
rect 61124 5964 68012 6020
rect 68068 5964 68078 6020
rect 93426 5964 93436 6020
rect 93492 5964 117628 6020
rect 117684 5964 117704 6020
rect 127586 5964 127596 6020
rect 127652 5964 139468 6020
rect 139524 5964 139534 6020
rect 194898 5964 194908 6020
rect 194964 5964 213164 6020
rect 213220 5964 213230 6020
rect 227602 5964 227612 6020
rect 227668 5964 255052 6020
rect 255108 5964 255118 6020
rect 267922 5964 267932 6020
rect 267988 5964 275996 6020
rect 276052 5964 276062 6020
rect 280578 5964 280588 6020
rect 280644 5964 344540 6020
rect 344596 5964 344606 6020
rect 364578 5964 364588 6020
rect 364644 5964 474012 6020
rect 474068 5964 474078 6020
rect 484642 5964 484652 6020
rect 484708 5964 508284 6020
rect 508340 5964 508350 6020
rect 13346 5852 13356 5908
rect 13412 5852 65548 5908
rect 65604 5852 65614 5908
rect 66770 5852 66780 5908
rect 66836 5852 83132 5908
rect 83188 5852 83198 5908
rect 87714 5852 87724 5908
rect 87780 5852 116172 5908
rect 116228 5852 116238 5908
rect 123890 5852 123900 5908
rect 123956 5852 125132 5908
rect 125188 5852 125198 5908
rect 125794 5852 125804 5908
rect 125860 5852 137900 5908
rect 137956 5852 137966 5908
rect 141026 5852 141036 5908
rect 141092 5852 147868 5908
rect 147924 5852 147934 5908
rect 179890 5852 179900 5908
rect 179956 5852 190316 5908
rect 190372 5852 190382 5908
rect 206658 5852 206668 5908
rect 206724 5852 230300 5908
rect 230356 5852 230366 5908
rect 233538 5852 233548 5908
rect 233604 5852 272188 5908
rect 272244 5852 272254 5908
rect 292338 5852 292348 5908
rect 292404 5852 363580 5908
rect 363636 5852 363646 5908
rect 409938 5852 409948 5908
rect 410004 5852 546364 5908
rect 546420 5852 546430 5908
rect 335122 5740 335132 5796
rect 335188 5740 338828 5796
rect 338884 5740 338894 5796
rect 17266 4956 17276 5012
rect 17332 4956 19292 5012
rect 19348 4956 19358 5012
rect 24882 4956 24892 5012
rect 24948 4956 27692 5012
rect 27748 4956 27758 5012
rect 40114 4956 40124 5012
rect 40180 4956 44492 5012
rect 44548 4956 44558 5012
rect 82898 4956 82908 5012
rect 82964 4956 90972 5012
rect 91028 4956 91038 5012
rect 133410 4956 133420 5012
rect 133476 4956 135212 5012
rect 135268 4956 135278 5012
rect 139122 4956 139132 5012
rect 139188 4956 140252 5012
rect 140308 4956 140318 5012
rect 146738 4956 146748 5012
rect 146804 4956 148652 5012
rect 148708 4956 148718 5012
rect 154354 4956 154364 5012
rect 154420 4956 156268 5012
rect 156324 4956 156334 5012
rect 158162 4956 158172 5012
rect 158228 4956 159628 5012
rect 159684 4956 159694 5012
rect 160066 4956 160076 5012
rect 160132 4956 161420 5012
rect 161476 4956 161486 5012
rect 166338 4956 166348 5012
rect 166404 4956 169372 5012
rect 169428 4956 169438 5012
rect 169698 4956 169708 5012
rect 169764 4956 173180 5012
rect 173236 4956 173246 5012
rect 180562 4956 180572 5012
rect 180628 4956 182700 5012
rect 182756 4956 182766 5012
rect 183138 4956 183148 5012
rect 183204 4956 194124 5012
rect 194180 4956 194190 5012
rect 215842 4956 215852 5012
rect 215908 4956 216972 5012
rect 217028 4956 217038 5012
rect 308242 4956 308252 5012
rect 308308 4956 310268 5012
rect 310324 4956 310334 5012
rect 373314 4956 373324 5012
rect 373380 4956 374780 5012
rect 374836 4956 374846 5012
rect 415762 4956 415772 5012
rect 415828 4956 416892 5012
rect 416948 4956 416958 5012
rect 456082 4956 456092 5012
rect 456148 4956 456988 5012
rect 457044 4956 457054 5012
rect 523282 4956 523292 5012
rect 523348 4956 525420 5012
rect 525476 4956 525486 5012
rect 560242 4956 560252 5012
rect 560308 4956 561596 5012
rect 561652 4956 561662 5012
rect 26786 4844 26796 4900
rect 26852 4844 34524 4900
rect 34580 4844 34590 4900
rect 68674 4844 68684 4900
rect 68740 4844 100940 4900
rect 100996 4844 101006 4900
rect 156146 4844 156156 4900
rect 156212 4844 157948 4900
rect 158004 4844 158014 4900
rect 169922 4844 169932 4900
rect 169988 4844 175084 4900
rect 175140 4844 175150 4900
rect 178882 4844 178892 4900
rect 178948 4844 184604 4900
rect 184660 4844 184670 4900
rect 188178 4844 188188 4900
rect 188244 4844 201740 4900
rect 201796 4844 201806 4900
rect 257058 4844 257068 4900
rect 257124 4844 308364 4900
rect 308420 4844 308430 4900
rect 62962 4732 62972 4788
rect 63028 4732 97468 4788
rect 97524 4732 97534 4788
rect 118178 4732 118188 4788
rect 118244 4732 132860 4788
rect 132916 4732 132926 4788
rect 193442 4732 193452 4788
rect 193508 4732 209356 4788
rect 209412 4732 209422 4788
rect 263778 4732 263788 4788
rect 263844 4732 319788 4788
rect 319844 4732 319854 4788
rect 404898 4732 404908 4788
rect 404964 4732 536844 4788
rect 536900 4732 536910 4788
rect 57250 4620 57260 4676
rect 57316 4620 94108 4676
rect 94164 4620 94184 4676
rect 101042 4620 101052 4676
rect 101108 4620 122668 4676
rect 122724 4620 122734 4676
rect 189858 4620 189868 4676
rect 189924 4620 205548 4676
rect 205604 4620 205614 4676
rect 223458 4620 223468 4676
rect 223524 4620 257068 4676
rect 257124 4620 257134 4676
rect 272290 4620 272300 4676
rect 272356 4620 331212 4676
rect 331268 4620 331278 4676
rect 408258 4620 408268 4676
rect 408324 4620 542668 4676
rect 542724 4620 542734 4676
rect 34402 4508 34412 4564
rect 34468 4508 36092 4564
rect 36148 4508 36158 4564
rect 51538 4508 51548 4564
rect 51604 4508 82908 4564
rect 82964 4508 82974 4564
rect 84028 4508 85708 4564
rect 85764 4508 85774 4564
rect 97234 4508 97244 4564
rect 97300 4508 119532 4564
rect 119588 4508 119598 4564
rect 174738 4508 174748 4564
rect 174804 4508 180796 4564
rect 180852 4508 180862 4564
rect 186498 4508 186508 4564
rect 186564 4508 199948 4564
rect 200004 4508 200014 4564
rect 201618 4508 201628 4564
rect 201684 4508 222684 4564
rect 222740 4508 222750 4564
rect 226818 4508 226828 4564
rect 226884 4508 262668 4564
rect 262724 4508 262734 4564
rect 275538 4508 275548 4564
rect 275604 4508 336924 4564
rect 336980 4508 336990 4564
rect 411618 4508 411628 4564
rect 411684 4508 548268 4564
rect 548324 4508 548334 4564
rect 84028 4452 84084 4508
rect 43922 4396 43932 4452
rect 43988 4396 84084 4452
rect 85810 4396 85820 4452
rect 85876 4396 112588 4452
rect 112644 4396 112654 4452
rect 114370 4396 114380 4452
rect 114436 4396 131068 4452
rect 131124 4396 131134 4452
rect 173058 4396 173068 4452
rect 173124 4396 178892 4452
rect 178948 4396 178958 4452
rect 188514 4396 188524 4452
rect 188580 4396 203644 4452
rect 203700 4396 203710 4452
rect 204978 4396 204988 4452
rect 205044 4396 228508 4452
rect 228564 4396 228574 4452
rect 230178 4396 230188 4452
rect 230244 4396 268380 4452
rect 268436 4396 268446 4452
rect 282258 4396 282268 4452
rect 282324 4396 348348 4452
rect 348404 4396 348414 4452
rect 420018 4396 420028 4452
rect 420084 4396 559692 4452
rect 559748 4396 559758 4452
rect 21074 4284 21084 4340
rect 21140 4284 70588 4340
rect 70644 4284 70664 4340
rect 80098 4284 80108 4340
rect 80164 4284 109452 4340
rect 109508 4284 109518 4340
rect 112466 4284 112476 4340
rect 112532 4284 129388 4340
rect 129444 4284 129454 4340
rect 150546 4284 150556 4340
rect 150612 4284 154588 4340
rect 154644 4284 154654 4340
rect 179778 4284 179788 4340
rect 179844 4284 188412 4340
rect 188468 4284 188478 4340
rect 191538 4284 191548 4340
rect 191604 4284 207452 4340
rect 207508 4284 207518 4340
rect 208338 4284 208348 4340
rect 208404 4284 234108 4340
rect 234164 4284 234174 4340
rect 245298 4284 245308 4340
rect 245364 4284 291228 4340
rect 291284 4284 291294 4340
rect 300738 4284 300748 4340
rect 300804 4284 376908 4340
rect 376964 4284 376974 4340
rect 423378 4284 423388 4340
rect 423444 4284 565404 4340
rect 565460 4284 565470 4340
rect 19170 4172 19180 4228
rect 19236 4172 68908 4228
rect 68964 4172 68974 4228
rect 74386 4172 74396 4228
rect 74452 4172 105868 4228
rect 105924 4172 105934 4228
rect 106754 4172 106764 4228
rect 106820 4172 126028 4228
rect 126084 4172 126094 4228
rect 135314 4172 135324 4228
rect 135380 4172 142716 4228
rect 142772 4172 142782 4228
rect 148642 4172 148652 4228
rect 148708 4172 152908 4228
rect 152964 4172 152974 4228
rect 178098 4172 178108 4228
rect 178164 4172 186508 4228
rect 186564 4172 186574 4228
rect 193218 4172 193228 4228
rect 193284 4172 211260 4228
rect 211316 4172 211326 4228
rect 211698 4172 211708 4228
rect 211764 4172 239820 4228
rect 239876 4172 239886 4228
rect 253698 4172 253708 4228
rect 253764 4172 302652 4228
rect 302708 4172 302718 4228
rect 304098 4172 304108 4228
rect 304164 4172 382620 4228
rect 382676 4172 382686 4228
rect 433458 4172 433468 4228
rect 433524 4172 584444 4228
rect 584500 4172 584510 4228
rect 131506 3836 131516 3892
rect 131572 3836 137788 3892
rect 137844 3836 137854 3892
rect 129602 3388 129612 3444
rect 129668 3388 132636 3444
rect 132692 3388 132702 3444
rect 339378 2604 339388 2660
rect 339444 2604 435932 2660
rect 435988 2604 435998 2660
rect 248658 2492 248668 2548
rect 248724 2492 295036 2548
rect 295092 2492 295102 2548
rect 376338 2492 376348 2548
rect 376404 2492 493052 2548
rect 493108 2492 493118 2548
<< via3 >>
rect 433468 439292 433524 439348
rect 433468 438508 433524 438564
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 6874 460350 7494 477922
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 6874 262350 7494 279922
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 6874 82350 7494 99922
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 6874 46350 7494 63922
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 6874 28350 7494 45922
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 6874 10350 7494 27922
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 508350 21774 525922
rect 21154 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 21774 508350
rect 21154 508226 21774 508294
rect 21154 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 21774 508226
rect 21154 508102 21774 508170
rect 21154 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 21774 508102
rect 21154 507978 21774 508046
rect 21154 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 21774 507978
rect 21154 490350 21774 507922
rect 21154 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 21774 490350
rect 21154 490226 21774 490294
rect 21154 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 21774 490226
rect 21154 490102 21774 490170
rect 21154 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 21774 490102
rect 21154 489978 21774 490046
rect 21154 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 21774 489978
rect 21154 472350 21774 489922
rect 21154 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 21774 472350
rect 21154 472226 21774 472294
rect 21154 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 21774 472226
rect 21154 472102 21774 472170
rect 21154 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 21774 472102
rect 21154 471978 21774 472046
rect 21154 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 21774 471978
rect 21154 454350 21774 471922
rect 21154 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 21774 454350
rect 21154 454226 21774 454294
rect 21154 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 21774 454226
rect 21154 454102 21774 454170
rect 21154 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 21774 454102
rect 21154 453978 21774 454046
rect 21154 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 21774 453978
rect 21154 436350 21774 453922
rect 21154 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 21774 436350
rect 21154 436226 21774 436294
rect 21154 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 21774 436226
rect 21154 436102 21774 436170
rect 21154 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 21774 436102
rect 21154 435978 21774 436046
rect 21154 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 21774 435978
rect 21154 418350 21774 435922
rect 21154 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 21774 418350
rect 21154 418226 21774 418294
rect 21154 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 21774 418226
rect 21154 418102 21774 418170
rect 21154 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 21774 418102
rect 21154 417978 21774 418046
rect 21154 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 21774 417978
rect 21154 400350 21774 417922
rect 21154 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 21774 400350
rect 21154 400226 21774 400294
rect 21154 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 21774 400226
rect 21154 400102 21774 400170
rect 21154 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 21774 400102
rect 21154 399978 21774 400046
rect 21154 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 21774 399978
rect 21154 382350 21774 399922
rect 21154 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 21774 382350
rect 21154 382226 21774 382294
rect 21154 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 21774 382226
rect 21154 382102 21774 382170
rect 21154 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 21774 382102
rect 21154 381978 21774 382046
rect 21154 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 21774 381978
rect 21154 364350 21774 381922
rect 21154 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 21774 364350
rect 21154 364226 21774 364294
rect 21154 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 21774 364226
rect 21154 364102 21774 364170
rect 21154 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 21774 364102
rect 21154 363978 21774 364046
rect 21154 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 21774 363978
rect 21154 346350 21774 363922
rect 21154 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 21774 346350
rect 21154 346226 21774 346294
rect 21154 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 21774 346226
rect 21154 346102 21774 346170
rect 21154 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 21774 346102
rect 21154 345978 21774 346046
rect 21154 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 21774 345978
rect 21154 328350 21774 345922
rect 21154 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 21774 328350
rect 21154 328226 21774 328294
rect 21154 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 21774 328226
rect 21154 328102 21774 328170
rect 21154 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 21774 328102
rect 21154 327978 21774 328046
rect 21154 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 21774 327978
rect 21154 310350 21774 327922
rect 21154 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 21774 310350
rect 21154 310226 21774 310294
rect 21154 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 21774 310226
rect 21154 310102 21774 310170
rect 21154 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 21774 310102
rect 21154 309978 21774 310046
rect 21154 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 21774 309978
rect 21154 292350 21774 309922
rect 21154 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 21774 292350
rect 21154 292226 21774 292294
rect 21154 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 21774 292226
rect 21154 292102 21774 292170
rect 21154 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 21774 292102
rect 21154 291978 21774 292046
rect 21154 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 21774 291978
rect 21154 274350 21774 291922
rect 21154 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 21774 274350
rect 21154 274226 21774 274294
rect 21154 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 21774 274226
rect 21154 274102 21774 274170
rect 21154 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 21774 274102
rect 21154 273978 21774 274046
rect 21154 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 21774 273978
rect 21154 256350 21774 273922
rect 21154 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 21774 256350
rect 21154 256226 21774 256294
rect 21154 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 21774 256226
rect 21154 256102 21774 256170
rect 21154 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 21774 256102
rect 21154 255978 21774 256046
rect 21154 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 21774 255978
rect 21154 238350 21774 255922
rect 21154 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 21774 238350
rect 21154 238226 21774 238294
rect 21154 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 21774 238226
rect 21154 238102 21774 238170
rect 21154 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 21774 238102
rect 21154 237978 21774 238046
rect 21154 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 21774 237978
rect 21154 220350 21774 237922
rect 21154 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 21774 220350
rect 21154 220226 21774 220294
rect 21154 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 21774 220226
rect 21154 220102 21774 220170
rect 21154 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 21774 220102
rect 21154 219978 21774 220046
rect 21154 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 21774 219978
rect 21154 202350 21774 219922
rect 21154 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 21774 202350
rect 21154 202226 21774 202294
rect 21154 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 21774 202226
rect 21154 202102 21774 202170
rect 21154 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 21774 202102
rect 21154 201978 21774 202046
rect 21154 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 21774 201978
rect 21154 184350 21774 201922
rect 21154 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 21774 184350
rect 21154 184226 21774 184294
rect 21154 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 21774 184226
rect 21154 184102 21774 184170
rect 21154 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 21774 184102
rect 21154 183978 21774 184046
rect 21154 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 21774 183978
rect 21154 166350 21774 183922
rect 21154 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 21774 166350
rect 21154 166226 21774 166294
rect 21154 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 21774 166226
rect 21154 166102 21774 166170
rect 21154 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 21774 166102
rect 21154 165978 21774 166046
rect 21154 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 21774 165978
rect 21154 148350 21774 165922
rect 21154 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 21774 148350
rect 21154 148226 21774 148294
rect 21154 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 21774 148226
rect 21154 148102 21774 148170
rect 21154 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 21774 148102
rect 21154 147978 21774 148046
rect 21154 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 21774 147978
rect 21154 130350 21774 147922
rect 21154 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 21774 130350
rect 21154 130226 21774 130294
rect 21154 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 21774 130226
rect 21154 130102 21774 130170
rect 21154 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 21774 130102
rect 21154 129978 21774 130046
rect 21154 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 21774 129978
rect 21154 112350 21774 129922
rect 21154 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 21774 112350
rect 21154 112226 21774 112294
rect 21154 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 21774 112226
rect 21154 112102 21774 112170
rect 21154 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 21774 112102
rect 21154 111978 21774 112046
rect 21154 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 21774 111978
rect 21154 94350 21774 111922
rect 21154 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 21774 94350
rect 21154 94226 21774 94294
rect 21154 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 21774 94226
rect 21154 94102 21774 94170
rect 21154 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 21774 94102
rect 21154 93978 21774 94046
rect 21154 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 21774 93978
rect 21154 76350 21774 93922
rect 21154 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 21774 76350
rect 21154 76226 21774 76294
rect 21154 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 21774 76226
rect 21154 76102 21774 76170
rect 21154 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 21774 76102
rect 21154 75978 21774 76046
rect 21154 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 21774 75978
rect 21154 58350 21774 75922
rect 21154 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 21774 58350
rect 21154 58226 21774 58294
rect 21154 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 21774 58226
rect 21154 58102 21774 58170
rect 21154 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 21774 58102
rect 21154 57978 21774 58046
rect 21154 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 21774 57978
rect 21154 40350 21774 57922
rect 21154 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 21774 40350
rect 21154 40226 21774 40294
rect 21154 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 21774 40226
rect 21154 40102 21774 40170
rect 21154 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 21774 40102
rect 21154 39978 21774 40046
rect 21154 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 21774 39978
rect 21154 22350 21774 39922
rect 21154 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 21774 22350
rect 21154 22226 21774 22294
rect 21154 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 21774 22226
rect 21154 22102 21774 22170
rect 21154 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 21774 22102
rect 21154 21978 21774 22046
rect 21154 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 21774 21978
rect 21154 4350 21774 21922
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 24874 514350 25494 531922
rect 24874 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 25494 514350
rect 24874 514226 25494 514294
rect 24874 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 25494 514226
rect 24874 514102 25494 514170
rect 24874 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 25494 514102
rect 24874 513978 25494 514046
rect 24874 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 25494 513978
rect 24874 496350 25494 513922
rect 24874 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 25494 496350
rect 24874 496226 25494 496294
rect 24874 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 25494 496226
rect 24874 496102 25494 496170
rect 24874 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 25494 496102
rect 24874 495978 25494 496046
rect 24874 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 25494 495978
rect 24874 478350 25494 495922
rect 24874 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 25494 478350
rect 24874 478226 25494 478294
rect 24874 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 25494 478226
rect 24874 478102 25494 478170
rect 24874 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 25494 478102
rect 24874 477978 25494 478046
rect 24874 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 25494 477978
rect 24874 460350 25494 477922
rect 24874 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 25494 460350
rect 24874 460226 25494 460294
rect 24874 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 25494 460226
rect 24874 460102 25494 460170
rect 24874 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 25494 460102
rect 24874 459978 25494 460046
rect 24874 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 25494 459978
rect 24874 442350 25494 459922
rect 24874 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 25494 442350
rect 24874 442226 25494 442294
rect 24874 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 25494 442226
rect 24874 442102 25494 442170
rect 24874 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 25494 442102
rect 24874 441978 25494 442046
rect 24874 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 25494 441978
rect 24874 424350 25494 441922
rect 24874 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 25494 424350
rect 24874 424226 25494 424294
rect 24874 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 25494 424226
rect 24874 424102 25494 424170
rect 24874 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 25494 424102
rect 24874 423978 25494 424046
rect 24874 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 25494 423978
rect 24874 406350 25494 423922
rect 24874 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 25494 406350
rect 24874 406226 25494 406294
rect 24874 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 25494 406226
rect 24874 406102 25494 406170
rect 24874 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 25494 406102
rect 24874 405978 25494 406046
rect 24874 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 25494 405978
rect 24874 388350 25494 405922
rect 24874 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 25494 388350
rect 24874 388226 25494 388294
rect 24874 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 25494 388226
rect 24874 388102 25494 388170
rect 24874 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 25494 388102
rect 24874 387978 25494 388046
rect 24874 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 25494 387978
rect 24874 370350 25494 387922
rect 24874 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 25494 370350
rect 24874 370226 25494 370294
rect 24874 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 25494 370226
rect 24874 370102 25494 370170
rect 24874 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 25494 370102
rect 24874 369978 25494 370046
rect 24874 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 25494 369978
rect 24874 352350 25494 369922
rect 24874 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 25494 352350
rect 24874 352226 25494 352294
rect 24874 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 25494 352226
rect 24874 352102 25494 352170
rect 24874 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 25494 352102
rect 24874 351978 25494 352046
rect 24874 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 25494 351978
rect 24874 334350 25494 351922
rect 24874 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 25494 334350
rect 24874 334226 25494 334294
rect 24874 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 25494 334226
rect 24874 334102 25494 334170
rect 24874 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 25494 334102
rect 24874 333978 25494 334046
rect 24874 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 25494 333978
rect 24874 316350 25494 333922
rect 24874 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 25494 316350
rect 24874 316226 25494 316294
rect 24874 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 25494 316226
rect 24874 316102 25494 316170
rect 24874 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 25494 316102
rect 24874 315978 25494 316046
rect 24874 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 25494 315978
rect 24874 298350 25494 315922
rect 24874 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 25494 298350
rect 24874 298226 25494 298294
rect 24874 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 25494 298226
rect 24874 298102 25494 298170
rect 24874 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 25494 298102
rect 24874 297978 25494 298046
rect 24874 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 25494 297978
rect 24874 280350 25494 297922
rect 24874 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 25494 280350
rect 24874 280226 25494 280294
rect 24874 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 25494 280226
rect 24874 280102 25494 280170
rect 24874 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 25494 280102
rect 24874 279978 25494 280046
rect 24874 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 25494 279978
rect 24874 262350 25494 279922
rect 24874 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 25494 262350
rect 24874 262226 25494 262294
rect 24874 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 25494 262226
rect 24874 262102 25494 262170
rect 24874 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 25494 262102
rect 24874 261978 25494 262046
rect 24874 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 25494 261978
rect 24874 244350 25494 261922
rect 24874 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 25494 244350
rect 24874 244226 25494 244294
rect 24874 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 25494 244226
rect 24874 244102 25494 244170
rect 24874 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 25494 244102
rect 24874 243978 25494 244046
rect 24874 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 25494 243978
rect 24874 226350 25494 243922
rect 24874 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 25494 226350
rect 24874 226226 25494 226294
rect 24874 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 25494 226226
rect 24874 226102 25494 226170
rect 24874 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 25494 226102
rect 24874 225978 25494 226046
rect 24874 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 25494 225978
rect 24874 208350 25494 225922
rect 24874 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 25494 208350
rect 24874 208226 25494 208294
rect 24874 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 25494 208226
rect 24874 208102 25494 208170
rect 24874 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 25494 208102
rect 24874 207978 25494 208046
rect 24874 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 25494 207978
rect 24874 190350 25494 207922
rect 24874 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 25494 190350
rect 24874 190226 25494 190294
rect 24874 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 25494 190226
rect 24874 190102 25494 190170
rect 24874 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 25494 190102
rect 24874 189978 25494 190046
rect 24874 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 25494 189978
rect 24874 172350 25494 189922
rect 24874 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 25494 172350
rect 24874 172226 25494 172294
rect 24874 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 25494 172226
rect 24874 172102 25494 172170
rect 24874 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 25494 172102
rect 24874 171978 25494 172046
rect 24874 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 25494 171978
rect 24874 154350 25494 171922
rect 24874 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 25494 154350
rect 24874 154226 25494 154294
rect 24874 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 25494 154226
rect 24874 154102 25494 154170
rect 24874 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 25494 154102
rect 24874 153978 25494 154046
rect 24874 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 25494 153978
rect 24874 136350 25494 153922
rect 24874 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 25494 136350
rect 24874 136226 25494 136294
rect 24874 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 25494 136226
rect 24874 136102 25494 136170
rect 24874 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 25494 136102
rect 24874 135978 25494 136046
rect 24874 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 25494 135978
rect 24874 118350 25494 135922
rect 24874 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 25494 118350
rect 24874 118226 25494 118294
rect 24874 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 25494 118226
rect 24874 118102 25494 118170
rect 24874 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 25494 118102
rect 24874 117978 25494 118046
rect 24874 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 25494 117978
rect 24874 100350 25494 117922
rect 24874 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 25494 100350
rect 24874 100226 25494 100294
rect 24874 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 25494 100226
rect 24874 100102 25494 100170
rect 24874 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 25494 100102
rect 24874 99978 25494 100046
rect 24874 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 25494 99978
rect 24874 82350 25494 99922
rect 24874 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 25494 82350
rect 24874 82226 25494 82294
rect 24874 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 25494 82226
rect 24874 82102 25494 82170
rect 24874 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 25494 82102
rect 24874 81978 25494 82046
rect 24874 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 25494 81978
rect 24874 64350 25494 81922
rect 24874 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 25494 64350
rect 24874 64226 25494 64294
rect 24874 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 25494 64226
rect 24874 64102 25494 64170
rect 24874 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 25494 64102
rect 24874 63978 25494 64046
rect 24874 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 25494 63978
rect 24874 46350 25494 63922
rect 24874 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 25494 46350
rect 24874 46226 25494 46294
rect 24874 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 25494 46226
rect 24874 46102 25494 46170
rect 24874 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 25494 46102
rect 24874 45978 25494 46046
rect 24874 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 25494 45978
rect 24874 28350 25494 45922
rect 24874 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 25494 28350
rect 24874 28226 25494 28294
rect 24874 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 25494 28226
rect 24874 28102 25494 28170
rect 24874 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 25494 28102
rect 24874 27978 25494 28046
rect 24874 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 25494 27978
rect 24874 10350 25494 27922
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 508350 39774 525922
rect 39154 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 39774 508350
rect 39154 508226 39774 508294
rect 39154 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 39774 508226
rect 39154 508102 39774 508170
rect 39154 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 39774 508102
rect 39154 507978 39774 508046
rect 39154 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 39774 507978
rect 39154 490350 39774 507922
rect 39154 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 39774 490350
rect 39154 490226 39774 490294
rect 39154 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 39774 490226
rect 39154 490102 39774 490170
rect 39154 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 39774 490102
rect 39154 489978 39774 490046
rect 39154 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 39774 489978
rect 39154 472350 39774 489922
rect 39154 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 39774 472350
rect 39154 472226 39774 472294
rect 39154 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 39774 472226
rect 39154 472102 39774 472170
rect 39154 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 39774 472102
rect 39154 471978 39774 472046
rect 39154 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 39774 471978
rect 39154 454350 39774 471922
rect 39154 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 39774 454350
rect 39154 454226 39774 454294
rect 39154 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 39774 454226
rect 39154 454102 39774 454170
rect 39154 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 39774 454102
rect 39154 453978 39774 454046
rect 39154 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 39774 453978
rect 39154 436350 39774 453922
rect 39154 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 39774 436350
rect 39154 436226 39774 436294
rect 39154 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 39774 436226
rect 39154 436102 39774 436170
rect 39154 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 39774 436102
rect 39154 435978 39774 436046
rect 39154 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 39774 435978
rect 39154 418350 39774 435922
rect 39154 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 39774 418350
rect 39154 418226 39774 418294
rect 39154 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 39774 418226
rect 39154 418102 39774 418170
rect 39154 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 39774 418102
rect 39154 417978 39774 418046
rect 39154 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 39774 417978
rect 39154 400350 39774 417922
rect 39154 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 39774 400350
rect 39154 400226 39774 400294
rect 39154 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 39774 400226
rect 39154 400102 39774 400170
rect 39154 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 39774 400102
rect 39154 399978 39774 400046
rect 39154 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 39774 399978
rect 39154 382350 39774 399922
rect 39154 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 39774 382350
rect 39154 382226 39774 382294
rect 39154 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 39774 382226
rect 39154 382102 39774 382170
rect 39154 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 39774 382102
rect 39154 381978 39774 382046
rect 39154 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 39774 381978
rect 39154 364350 39774 381922
rect 39154 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 39774 364350
rect 39154 364226 39774 364294
rect 39154 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 39774 364226
rect 39154 364102 39774 364170
rect 39154 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 39774 364102
rect 39154 363978 39774 364046
rect 39154 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 39774 363978
rect 39154 346350 39774 363922
rect 39154 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 39774 346350
rect 39154 346226 39774 346294
rect 39154 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 39774 346226
rect 39154 346102 39774 346170
rect 39154 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 39774 346102
rect 39154 345978 39774 346046
rect 39154 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 39774 345978
rect 39154 328350 39774 345922
rect 39154 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 39774 328350
rect 39154 328226 39774 328294
rect 39154 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 39774 328226
rect 39154 328102 39774 328170
rect 39154 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 39774 328102
rect 39154 327978 39774 328046
rect 39154 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 39774 327978
rect 39154 310350 39774 327922
rect 39154 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 39774 310350
rect 39154 310226 39774 310294
rect 39154 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 39774 310226
rect 39154 310102 39774 310170
rect 39154 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 39774 310102
rect 39154 309978 39774 310046
rect 39154 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 39774 309978
rect 39154 292350 39774 309922
rect 39154 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 39774 292350
rect 39154 292226 39774 292294
rect 39154 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 39774 292226
rect 39154 292102 39774 292170
rect 39154 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 39774 292102
rect 39154 291978 39774 292046
rect 39154 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 39774 291978
rect 39154 274350 39774 291922
rect 39154 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 39774 274350
rect 39154 274226 39774 274294
rect 39154 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 39774 274226
rect 39154 274102 39774 274170
rect 39154 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 39774 274102
rect 39154 273978 39774 274046
rect 39154 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 39774 273978
rect 39154 256350 39774 273922
rect 39154 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 39774 256350
rect 39154 256226 39774 256294
rect 39154 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 39774 256226
rect 39154 256102 39774 256170
rect 39154 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 39774 256102
rect 39154 255978 39774 256046
rect 39154 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 39774 255978
rect 39154 238350 39774 255922
rect 39154 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 39774 238350
rect 39154 238226 39774 238294
rect 39154 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 39774 238226
rect 39154 238102 39774 238170
rect 39154 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 39774 238102
rect 39154 237978 39774 238046
rect 39154 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 39774 237978
rect 39154 220350 39774 237922
rect 39154 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 39774 220350
rect 39154 220226 39774 220294
rect 39154 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 39774 220226
rect 39154 220102 39774 220170
rect 39154 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 39774 220102
rect 39154 219978 39774 220046
rect 39154 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 39774 219978
rect 39154 202350 39774 219922
rect 39154 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 39774 202350
rect 39154 202226 39774 202294
rect 39154 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 39774 202226
rect 39154 202102 39774 202170
rect 39154 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 39774 202102
rect 39154 201978 39774 202046
rect 39154 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 39774 201978
rect 39154 184350 39774 201922
rect 39154 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 39774 184350
rect 39154 184226 39774 184294
rect 39154 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 39774 184226
rect 39154 184102 39774 184170
rect 39154 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 39774 184102
rect 39154 183978 39774 184046
rect 39154 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 39774 183978
rect 39154 166350 39774 183922
rect 39154 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 39774 166350
rect 39154 166226 39774 166294
rect 39154 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 39774 166226
rect 39154 166102 39774 166170
rect 39154 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 39774 166102
rect 39154 165978 39774 166046
rect 39154 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 39774 165978
rect 39154 148350 39774 165922
rect 39154 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 39774 148350
rect 39154 148226 39774 148294
rect 39154 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 39774 148226
rect 39154 148102 39774 148170
rect 39154 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 39774 148102
rect 39154 147978 39774 148046
rect 39154 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 39774 147978
rect 39154 130350 39774 147922
rect 39154 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 39774 130350
rect 39154 130226 39774 130294
rect 39154 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 39774 130226
rect 39154 130102 39774 130170
rect 39154 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 39774 130102
rect 39154 129978 39774 130046
rect 39154 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 39774 129978
rect 39154 112350 39774 129922
rect 39154 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 39774 112350
rect 39154 112226 39774 112294
rect 39154 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 39774 112226
rect 39154 112102 39774 112170
rect 39154 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 39774 112102
rect 39154 111978 39774 112046
rect 39154 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 39774 111978
rect 39154 94350 39774 111922
rect 39154 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 39774 94350
rect 39154 94226 39774 94294
rect 39154 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 39774 94226
rect 39154 94102 39774 94170
rect 39154 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 39774 94102
rect 39154 93978 39774 94046
rect 39154 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 39774 93978
rect 39154 76350 39774 93922
rect 39154 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 39774 76350
rect 39154 76226 39774 76294
rect 39154 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 39774 76226
rect 39154 76102 39774 76170
rect 39154 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 39774 76102
rect 39154 75978 39774 76046
rect 39154 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 39774 75978
rect 39154 58350 39774 75922
rect 39154 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 39774 58350
rect 39154 58226 39774 58294
rect 39154 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 39774 58226
rect 39154 58102 39774 58170
rect 39154 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 39774 58102
rect 39154 57978 39774 58046
rect 39154 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 39774 57978
rect 39154 40350 39774 57922
rect 39154 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 39774 40350
rect 39154 40226 39774 40294
rect 39154 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 39774 40226
rect 39154 40102 39774 40170
rect 39154 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 39774 40102
rect 39154 39978 39774 40046
rect 39154 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 39774 39978
rect 39154 22350 39774 39922
rect 39154 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 39774 22350
rect 39154 22226 39774 22294
rect 39154 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 39774 22226
rect 39154 22102 39774 22170
rect 39154 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 39774 22102
rect 39154 21978 39774 22046
rect 39154 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 39774 21978
rect 39154 4350 39774 21922
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 514350 43494 531922
rect 42874 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 43494 514350
rect 42874 514226 43494 514294
rect 42874 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 43494 514226
rect 42874 514102 43494 514170
rect 42874 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 43494 514102
rect 42874 513978 43494 514046
rect 42874 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 43494 513978
rect 42874 496350 43494 513922
rect 42874 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 43494 496350
rect 42874 496226 43494 496294
rect 42874 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 43494 496226
rect 42874 496102 43494 496170
rect 42874 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 43494 496102
rect 42874 495978 43494 496046
rect 42874 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 43494 495978
rect 42874 478350 43494 495922
rect 42874 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 43494 478350
rect 42874 478226 43494 478294
rect 42874 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 43494 478226
rect 42874 478102 43494 478170
rect 42874 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 43494 478102
rect 42874 477978 43494 478046
rect 42874 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 43494 477978
rect 42874 460350 43494 477922
rect 42874 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 43494 460350
rect 42874 460226 43494 460294
rect 42874 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 43494 460226
rect 42874 460102 43494 460170
rect 42874 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 43494 460102
rect 42874 459978 43494 460046
rect 42874 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 43494 459978
rect 42874 442350 43494 459922
rect 42874 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 43494 442350
rect 42874 442226 43494 442294
rect 42874 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 43494 442226
rect 42874 442102 43494 442170
rect 42874 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 43494 442102
rect 42874 441978 43494 442046
rect 42874 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 43494 441978
rect 42874 424350 43494 441922
rect 42874 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 43494 424350
rect 42874 424226 43494 424294
rect 42874 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 43494 424226
rect 42874 424102 43494 424170
rect 42874 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 43494 424102
rect 42874 423978 43494 424046
rect 42874 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 43494 423978
rect 42874 406350 43494 423922
rect 42874 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 43494 406350
rect 42874 406226 43494 406294
rect 42874 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 43494 406226
rect 42874 406102 43494 406170
rect 42874 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 43494 406102
rect 42874 405978 43494 406046
rect 42874 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 43494 405978
rect 42874 388350 43494 405922
rect 42874 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 43494 388350
rect 42874 388226 43494 388294
rect 42874 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 43494 388226
rect 42874 388102 43494 388170
rect 42874 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 43494 388102
rect 42874 387978 43494 388046
rect 42874 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 43494 387978
rect 42874 370350 43494 387922
rect 42874 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 43494 370350
rect 42874 370226 43494 370294
rect 42874 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 43494 370226
rect 42874 370102 43494 370170
rect 42874 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 43494 370102
rect 42874 369978 43494 370046
rect 42874 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 43494 369978
rect 42874 352350 43494 369922
rect 42874 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 43494 352350
rect 42874 352226 43494 352294
rect 42874 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 43494 352226
rect 42874 352102 43494 352170
rect 42874 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 43494 352102
rect 42874 351978 43494 352046
rect 42874 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 43494 351978
rect 42874 334350 43494 351922
rect 42874 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 43494 334350
rect 42874 334226 43494 334294
rect 42874 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 43494 334226
rect 42874 334102 43494 334170
rect 42874 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 43494 334102
rect 42874 333978 43494 334046
rect 42874 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 43494 333978
rect 42874 316350 43494 333922
rect 42874 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 43494 316350
rect 42874 316226 43494 316294
rect 42874 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 43494 316226
rect 42874 316102 43494 316170
rect 42874 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 43494 316102
rect 42874 315978 43494 316046
rect 42874 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 43494 315978
rect 42874 298350 43494 315922
rect 42874 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 43494 298350
rect 42874 298226 43494 298294
rect 42874 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 43494 298226
rect 42874 298102 43494 298170
rect 42874 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 43494 298102
rect 42874 297978 43494 298046
rect 42874 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 43494 297978
rect 42874 280350 43494 297922
rect 42874 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 43494 280350
rect 42874 280226 43494 280294
rect 42874 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 43494 280226
rect 42874 280102 43494 280170
rect 42874 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 43494 280102
rect 42874 279978 43494 280046
rect 42874 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 43494 279978
rect 42874 262350 43494 279922
rect 42874 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 43494 262350
rect 42874 262226 43494 262294
rect 42874 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 43494 262226
rect 42874 262102 43494 262170
rect 42874 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 43494 262102
rect 42874 261978 43494 262046
rect 42874 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 43494 261978
rect 42874 244350 43494 261922
rect 42874 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 43494 244350
rect 42874 244226 43494 244294
rect 42874 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 43494 244226
rect 42874 244102 43494 244170
rect 42874 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 43494 244102
rect 42874 243978 43494 244046
rect 42874 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 43494 243978
rect 42874 226350 43494 243922
rect 42874 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 43494 226350
rect 42874 226226 43494 226294
rect 42874 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 43494 226226
rect 42874 226102 43494 226170
rect 42874 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 43494 226102
rect 42874 225978 43494 226046
rect 42874 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 43494 225978
rect 42874 208350 43494 225922
rect 42874 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 43494 208350
rect 42874 208226 43494 208294
rect 42874 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 43494 208226
rect 42874 208102 43494 208170
rect 42874 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 43494 208102
rect 42874 207978 43494 208046
rect 42874 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 43494 207978
rect 42874 190350 43494 207922
rect 42874 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 43494 190350
rect 42874 190226 43494 190294
rect 42874 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 43494 190226
rect 42874 190102 43494 190170
rect 42874 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 43494 190102
rect 42874 189978 43494 190046
rect 42874 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 43494 189978
rect 42874 172350 43494 189922
rect 42874 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 43494 172350
rect 42874 172226 43494 172294
rect 42874 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 43494 172226
rect 42874 172102 43494 172170
rect 42874 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 43494 172102
rect 42874 171978 43494 172046
rect 42874 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 43494 171978
rect 42874 154350 43494 171922
rect 42874 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 43494 154350
rect 42874 154226 43494 154294
rect 42874 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 43494 154226
rect 42874 154102 43494 154170
rect 42874 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 43494 154102
rect 42874 153978 43494 154046
rect 42874 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 43494 153978
rect 42874 136350 43494 153922
rect 42874 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 43494 136350
rect 42874 136226 43494 136294
rect 42874 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 43494 136226
rect 42874 136102 43494 136170
rect 42874 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 43494 136102
rect 42874 135978 43494 136046
rect 42874 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 43494 135978
rect 42874 118350 43494 135922
rect 42874 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 43494 118350
rect 42874 118226 43494 118294
rect 42874 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 43494 118226
rect 42874 118102 43494 118170
rect 42874 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 43494 118102
rect 42874 117978 43494 118046
rect 42874 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 43494 117978
rect 42874 100350 43494 117922
rect 42874 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 43494 100350
rect 42874 100226 43494 100294
rect 42874 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 43494 100226
rect 42874 100102 43494 100170
rect 42874 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 43494 100102
rect 42874 99978 43494 100046
rect 42874 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 43494 99978
rect 42874 82350 43494 99922
rect 42874 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 43494 82350
rect 42874 82226 43494 82294
rect 42874 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 43494 82226
rect 42874 82102 43494 82170
rect 42874 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 43494 82102
rect 42874 81978 43494 82046
rect 42874 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 43494 81978
rect 42874 64350 43494 81922
rect 42874 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 43494 64350
rect 42874 64226 43494 64294
rect 42874 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 43494 64226
rect 42874 64102 43494 64170
rect 42874 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 43494 64102
rect 42874 63978 43494 64046
rect 42874 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 43494 63978
rect 42874 46350 43494 63922
rect 42874 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 43494 46350
rect 42874 46226 43494 46294
rect 42874 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 43494 46226
rect 42874 46102 43494 46170
rect 42874 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 43494 46102
rect 42874 45978 43494 46046
rect 42874 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 43494 45978
rect 42874 28350 43494 45922
rect 42874 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 43494 28350
rect 42874 28226 43494 28294
rect 42874 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 43494 28226
rect 42874 28102 43494 28170
rect 42874 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 43494 28102
rect 42874 27978 43494 28046
rect 42874 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 43494 27978
rect 42874 10350 43494 27922
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 57154 508350 57774 525922
rect 57154 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 57774 508350
rect 57154 508226 57774 508294
rect 57154 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 57774 508226
rect 57154 508102 57774 508170
rect 57154 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 57774 508102
rect 57154 507978 57774 508046
rect 57154 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 57774 507978
rect 57154 490350 57774 507922
rect 57154 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 57774 490350
rect 57154 490226 57774 490294
rect 57154 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 57774 490226
rect 57154 490102 57774 490170
rect 57154 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 57774 490102
rect 57154 489978 57774 490046
rect 57154 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 57774 489978
rect 57154 472350 57774 489922
rect 57154 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 57774 472350
rect 57154 472226 57774 472294
rect 57154 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 57774 472226
rect 57154 472102 57774 472170
rect 57154 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 57774 472102
rect 57154 471978 57774 472046
rect 57154 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 57774 471978
rect 57154 454350 57774 471922
rect 57154 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 57774 454350
rect 57154 454226 57774 454294
rect 57154 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 57774 454226
rect 57154 454102 57774 454170
rect 57154 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 57774 454102
rect 57154 453978 57774 454046
rect 57154 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 57774 453978
rect 57154 436350 57774 453922
rect 57154 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 57774 436350
rect 57154 436226 57774 436294
rect 57154 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 57774 436226
rect 57154 436102 57774 436170
rect 57154 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 57774 436102
rect 57154 435978 57774 436046
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 514350 61494 531922
rect 60874 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 61494 514350
rect 60874 514226 61494 514294
rect 60874 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 61494 514226
rect 60874 514102 61494 514170
rect 60874 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 61494 514102
rect 60874 513978 61494 514046
rect 60874 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 61494 513978
rect 60874 496350 61494 513922
rect 60874 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 61494 496350
rect 60874 496226 61494 496294
rect 60874 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 61494 496226
rect 60874 496102 61494 496170
rect 60874 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 61494 496102
rect 60874 495978 61494 496046
rect 60874 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 61494 495978
rect 60874 478350 61494 495922
rect 60874 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 61494 478350
rect 60874 478226 61494 478294
rect 60874 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 61494 478226
rect 60874 478102 61494 478170
rect 60874 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 61494 478102
rect 60874 477978 61494 478046
rect 60874 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 61494 477978
rect 60874 460350 61494 477922
rect 60874 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 61494 460350
rect 60874 460226 61494 460294
rect 60874 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 61494 460226
rect 60874 460102 61494 460170
rect 60874 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 61494 460102
rect 60874 459978 61494 460046
rect 60874 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 61494 459978
rect 60874 442350 61494 459922
rect 60874 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 61494 442350
rect 60874 442226 61494 442294
rect 60874 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 61494 442226
rect 60874 442102 61494 442170
rect 60874 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 61494 442102
rect 60874 441978 61494 442046
rect 60874 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 61494 441978
rect 60874 436006 61494 441922
rect 75154 597212 75774 598268
rect 75154 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 75774 597212
rect 75154 597088 75774 597156
rect 75154 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 75774 597088
rect 75154 596964 75774 597032
rect 75154 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 75774 596964
rect 75154 596840 75774 596908
rect 75154 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 75774 596840
rect 75154 580350 75774 596784
rect 75154 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 75774 580350
rect 75154 580226 75774 580294
rect 75154 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 75774 580226
rect 75154 580102 75774 580170
rect 75154 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 75774 580102
rect 75154 579978 75774 580046
rect 75154 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 75774 579978
rect 75154 562350 75774 579922
rect 75154 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 75774 562350
rect 75154 562226 75774 562294
rect 75154 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 75774 562226
rect 75154 562102 75774 562170
rect 75154 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 75774 562102
rect 75154 561978 75774 562046
rect 75154 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 75774 561978
rect 75154 544350 75774 561922
rect 75154 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 75774 544350
rect 75154 544226 75774 544294
rect 75154 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 75774 544226
rect 75154 544102 75774 544170
rect 75154 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 75774 544102
rect 75154 543978 75774 544046
rect 75154 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 75774 543978
rect 75154 526350 75774 543922
rect 75154 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 75774 526350
rect 75154 526226 75774 526294
rect 75154 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 75774 526226
rect 75154 526102 75774 526170
rect 75154 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 75774 526102
rect 75154 525978 75774 526046
rect 75154 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 75774 525978
rect 75154 508350 75774 525922
rect 75154 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 75774 508350
rect 75154 508226 75774 508294
rect 75154 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 75774 508226
rect 75154 508102 75774 508170
rect 75154 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 75774 508102
rect 75154 507978 75774 508046
rect 75154 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 75774 507978
rect 75154 490350 75774 507922
rect 75154 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 75774 490350
rect 75154 490226 75774 490294
rect 75154 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 75774 490226
rect 75154 490102 75774 490170
rect 75154 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 75774 490102
rect 75154 489978 75774 490046
rect 75154 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 75774 489978
rect 75154 472350 75774 489922
rect 75154 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 75774 472350
rect 75154 472226 75774 472294
rect 75154 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 75774 472226
rect 75154 472102 75774 472170
rect 75154 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 75774 472102
rect 75154 471978 75774 472046
rect 75154 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 75774 471978
rect 75154 454350 75774 471922
rect 75154 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 75774 454350
rect 75154 454226 75774 454294
rect 75154 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 75774 454226
rect 75154 454102 75774 454170
rect 75154 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 75774 454102
rect 75154 453978 75774 454046
rect 75154 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 75774 453978
rect 64448 436317 64768 436380
rect 64448 436261 64518 436317
rect 64574 436261 64642 436317
rect 64698 436261 64768 436317
rect 64448 436193 64768 436261
rect 64448 436137 64518 436193
rect 64574 436137 64642 436193
rect 64698 436137 64768 436193
rect 64448 436069 64768 436137
rect 64448 436013 64518 436069
rect 64574 436013 64642 436069
rect 64698 436013 64768 436069
rect 57154 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 57774 435978
rect 57154 418350 57774 435922
rect 64448 435945 64768 436013
rect 75154 436378 75774 453922
rect 75154 436322 75250 436378
rect 75306 436322 75374 436378
rect 75430 436322 75498 436378
rect 75554 436322 75622 436378
rect 75678 436322 75774 436378
rect 75154 436254 75774 436322
rect 75154 436198 75250 436254
rect 75306 436198 75374 436254
rect 75430 436198 75498 436254
rect 75554 436198 75622 436254
rect 75678 436198 75774 436254
rect 75154 436130 75774 436198
rect 75154 436074 75250 436130
rect 75306 436074 75374 436130
rect 75430 436074 75498 436130
rect 75554 436074 75622 436130
rect 75678 436074 75774 436130
rect 75154 436006 75774 436074
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 514350 79494 531922
rect 78874 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 79494 514350
rect 78874 514226 79494 514294
rect 78874 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 79494 514226
rect 78874 514102 79494 514170
rect 78874 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 79494 514102
rect 78874 513978 79494 514046
rect 78874 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 79494 513978
rect 78874 496350 79494 513922
rect 78874 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 79494 496350
rect 78874 496226 79494 496294
rect 78874 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 79494 496226
rect 78874 496102 79494 496170
rect 78874 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 79494 496102
rect 78874 495978 79494 496046
rect 78874 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 79494 495978
rect 78874 478350 79494 495922
rect 78874 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 79494 478350
rect 78874 478226 79494 478294
rect 78874 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 79494 478226
rect 78874 478102 79494 478170
rect 78874 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 79494 478102
rect 78874 477978 79494 478046
rect 78874 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 79494 477978
rect 78874 460350 79494 477922
rect 78874 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 79494 460350
rect 78874 460226 79494 460294
rect 78874 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 79494 460226
rect 78874 460102 79494 460170
rect 78874 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 79494 460102
rect 78874 459978 79494 460046
rect 78874 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 79494 459978
rect 78874 442350 79494 459922
rect 78874 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 79494 442350
rect 78874 442226 79494 442294
rect 78874 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 79494 442226
rect 78874 442102 79494 442170
rect 78874 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 79494 442102
rect 78874 441978 79494 442046
rect 78874 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 79494 441978
rect 78874 436006 79494 441922
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 93154 508350 93774 525922
rect 93154 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 93774 508350
rect 93154 508226 93774 508294
rect 93154 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 93774 508226
rect 93154 508102 93774 508170
rect 93154 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 93774 508102
rect 93154 507978 93774 508046
rect 93154 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 93774 507978
rect 93154 490350 93774 507922
rect 93154 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 93774 490350
rect 93154 490226 93774 490294
rect 93154 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 93774 490226
rect 93154 490102 93774 490170
rect 93154 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 93774 490102
rect 93154 489978 93774 490046
rect 93154 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 93774 489978
rect 93154 472350 93774 489922
rect 93154 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 93774 472350
rect 93154 472226 93774 472294
rect 93154 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 93774 472226
rect 93154 472102 93774 472170
rect 93154 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 93774 472102
rect 93154 471978 93774 472046
rect 93154 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 93774 471978
rect 93154 454350 93774 471922
rect 93154 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 93774 454350
rect 93154 454226 93774 454294
rect 93154 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 93774 454226
rect 93154 454102 93774 454170
rect 93154 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 93774 454102
rect 93154 453978 93774 454046
rect 93154 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 93774 453978
rect 93154 436378 93774 453922
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 514350 97494 531922
rect 96874 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 97494 514350
rect 96874 514226 97494 514294
rect 96874 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 97494 514226
rect 96874 514102 97494 514170
rect 96874 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 97494 514102
rect 96874 513978 97494 514046
rect 96874 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 97494 513978
rect 96874 496350 97494 513922
rect 96874 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 97494 496350
rect 96874 496226 97494 496294
rect 96874 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 97494 496226
rect 96874 496102 97494 496170
rect 96874 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 97494 496102
rect 96874 495978 97494 496046
rect 96874 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 97494 495978
rect 96874 478350 97494 495922
rect 96874 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 97494 478350
rect 96874 478226 97494 478294
rect 96874 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 97494 478226
rect 96874 478102 97494 478170
rect 96874 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 97494 478102
rect 96874 477978 97494 478046
rect 96874 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 97494 477978
rect 96874 460350 97494 477922
rect 96874 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 97494 460350
rect 96874 460226 97494 460294
rect 96874 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 97494 460226
rect 96874 460102 97494 460170
rect 96874 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 97494 460102
rect 96874 459978 97494 460046
rect 96874 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 97494 459978
rect 96874 442350 97494 459922
rect 96874 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 97494 442350
rect 96874 442226 97494 442294
rect 96874 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 97494 442226
rect 96874 442102 97494 442170
rect 96874 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 97494 442102
rect 96874 441978 97494 442046
rect 96874 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 97494 441978
rect 93154 436322 93250 436378
rect 93306 436322 93374 436378
rect 93430 436322 93498 436378
rect 93554 436322 93622 436378
rect 93678 436322 93774 436378
rect 93154 436254 93774 436322
rect 93154 436198 93250 436254
rect 93306 436198 93374 436254
rect 93430 436198 93498 436254
rect 93554 436198 93622 436254
rect 93678 436198 93774 436254
rect 93154 436130 93774 436198
rect 93154 436074 93250 436130
rect 93306 436074 93374 436130
rect 93430 436074 93498 436130
rect 93554 436074 93622 436130
rect 93678 436074 93774 436130
rect 93154 436006 93774 436074
rect 95168 436317 95488 436380
rect 95168 436261 95238 436317
rect 95294 436261 95362 436317
rect 95418 436261 95488 436317
rect 95168 436193 95488 436261
rect 95168 436137 95238 436193
rect 95294 436137 95362 436193
rect 95418 436137 95488 436193
rect 95168 436069 95488 436137
rect 95168 436013 95238 436069
rect 95294 436013 95362 436069
rect 95418 436013 95488 436069
rect 64448 435889 64518 435945
rect 64574 435889 64642 435945
rect 64698 435889 64768 435945
rect 64448 435826 64768 435889
rect 95168 435945 95488 436013
rect 96874 436006 97494 441922
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 111154 508350 111774 525922
rect 111154 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 111774 508350
rect 111154 508226 111774 508294
rect 111154 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 111774 508226
rect 111154 508102 111774 508170
rect 111154 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 111774 508102
rect 111154 507978 111774 508046
rect 111154 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 111774 507978
rect 111154 490350 111774 507922
rect 111154 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 111774 490350
rect 111154 490226 111774 490294
rect 111154 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 111774 490226
rect 111154 490102 111774 490170
rect 111154 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 111774 490102
rect 111154 489978 111774 490046
rect 111154 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 111774 489978
rect 111154 472350 111774 489922
rect 111154 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 111774 472350
rect 111154 472226 111774 472294
rect 111154 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 111774 472226
rect 111154 472102 111774 472170
rect 111154 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 111774 472102
rect 111154 471978 111774 472046
rect 111154 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 111774 471978
rect 111154 454350 111774 471922
rect 111154 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 111774 454350
rect 111154 454226 111774 454294
rect 111154 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 111774 454226
rect 111154 454102 111774 454170
rect 111154 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 111774 454102
rect 111154 453978 111774 454046
rect 111154 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 111774 453978
rect 111154 436378 111774 453922
rect 111154 436322 111250 436378
rect 111306 436322 111374 436378
rect 111430 436322 111498 436378
rect 111554 436322 111622 436378
rect 111678 436322 111774 436378
rect 111154 436254 111774 436322
rect 111154 436198 111250 436254
rect 111306 436198 111374 436254
rect 111430 436198 111498 436254
rect 111554 436198 111622 436254
rect 111678 436198 111774 436254
rect 111154 436130 111774 436198
rect 111154 436074 111250 436130
rect 111306 436074 111374 436130
rect 111430 436074 111498 436130
rect 111554 436074 111622 436130
rect 111678 436074 111774 436130
rect 111154 436006 111774 436074
rect 114874 598172 115494 598268
rect 114874 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 115494 598172
rect 114874 598048 115494 598116
rect 114874 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 115494 598048
rect 114874 597924 115494 597992
rect 114874 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 115494 597924
rect 114874 597800 115494 597868
rect 114874 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 115494 597800
rect 114874 586350 115494 597744
rect 114874 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 115494 586350
rect 114874 586226 115494 586294
rect 114874 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 115494 586226
rect 114874 586102 115494 586170
rect 114874 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 115494 586102
rect 114874 585978 115494 586046
rect 114874 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 115494 585978
rect 114874 568350 115494 585922
rect 114874 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 115494 568350
rect 114874 568226 115494 568294
rect 114874 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 115494 568226
rect 114874 568102 115494 568170
rect 114874 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 115494 568102
rect 114874 567978 115494 568046
rect 114874 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 115494 567978
rect 114874 550350 115494 567922
rect 114874 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 115494 550350
rect 114874 550226 115494 550294
rect 114874 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 115494 550226
rect 114874 550102 115494 550170
rect 114874 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 115494 550102
rect 114874 549978 115494 550046
rect 114874 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 115494 549978
rect 114874 532350 115494 549922
rect 114874 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 115494 532350
rect 114874 532226 115494 532294
rect 114874 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 115494 532226
rect 114874 532102 115494 532170
rect 114874 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 115494 532102
rect 114874 531978 115494 532046
rect 114874 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 115494 531978
rect 114874 514350 115494 531922
rect 114874 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 115494 514350
rect 114874 514226 115494 514294
rect 114874 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 115494 514226
rect 114874 514102 115494 514170
rect 114874 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 115494 514102
rect 114874 513978 115494 514046
rect 114874 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 115494 513978
rect 114874 496350 115494 513922
rect 114874 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 115494 496350
rect 114874 496226 115494 496294
rect 114874 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 115494 496226
rect 114874 496102 115494 496170
rect 114874 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 115494 496102
rect 114874 495978 115494 496046
rect 114874 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 115494 495978
rect 114874 478350 115494 495922
rect 114874 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 115494 478350
rect 114874 478226 115494 478294
rect 114874 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 115494 478226
rect 114874 478102 115494 478170
rect 114874 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 115494 478102
rect 114874 477978 115494 478046
rect 114874 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 115494 477978
rect 114874 460350 115494 477922
rect 114874 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 115494 460350
rect 114874 460226 115494 460294
rect 114874 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 115494 460226
rect 114874 460102 115494 460170
rect 114874 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 115494 460102
rect 114874 459978 115494 460046
rect 114874 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 115494 459978
rect 114874 442350 115494 459922
rect 114874 442294 114970 442350
rect 115026 442294 115094 442350
rect 115150 442294 115218 442350
rect 115274 442294 115342 442350
rect 115398 442294 115494 442350
rect 114874 442226 115494 442294
rect 114874 442170 114970 442226
rect 115026 442170 115094 442226
rect 115150 442170 115218 442226
rect 115274 442170 115342 442226
rect 115398 442170 115494 442226
rect 114874 442102 115494 442170
rect 114874 442046 114970 442102
rect 115026 442046 115094 442102
rect 115150 442046 115218 442102
rect 115274 442046 115342 442102
rect 115398 442046 115494 442102
rect 114874 441978 115494 442046
rect 114874 441922 114970 441978
rect 115026 441922 115094 441978
rect 115150 441922 115218 441978
rect 115274 441922 115342 441978
rect 115398 441922 115494 441978
rect 114874 436006 115494 441922
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 526350 129774 543922
rect 129154 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 129774 526350
rect 129154 526226 129774 526294
rect 129154 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 129774 526226
rect 129154 526102 129774 526170
rect 129154 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 129774 526102
rect 129154 525978 129774 526046
rect 129154 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 129774 525978
rect 129154 508350 129774 525922
rect 129154 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 129774 508350
rect 129154 508226 129774 508294
rect 129154 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 129774 508226
rect 129154 508102 129774 508170
rect 129154 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 129774 508102
rect 129154 507978 129774 508046
rect 129154 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 129774 507978
rect 129154 490350 129774 507922
rect 129154 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 129774 490350
rect 129154 490226 129774 490294
rect 129154 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 129774 490226
rect 129154 490102 129774 490170
rect 129154 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 129774 490102
rect 129154 489978 129774 490046
rect 129154 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 129774 489978
rect 129154 472350 129774 489922
rect 129154 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 129774 472350
rect 129154 472226 129774 472294
rect 129154 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 129774 472226
rect 129154 472102 129774 472170
rect 129154 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 129774 472102
rect 129154 471978 129774 472046
rect 129154 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 129774 471978
rect 129154 454350 129774 471922
rect 129154 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 129774 454350
rect 129154 454226 129774 454294
rect 129154 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 129774 454226
rect 129154 454102 129774 454170
rect 129154 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 129774 454102
rect 129154 453978 129774 454046
rect 129154 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 129774 453978
rect 125888 436317 126208 436380
rect 125888 436261 125958 436317
rect 126014 436261 126082 436317
rect 126138 436261 126208 436317
rect 125888 436193 126208 436261
rect 125888 436137 125958 436193
rect 126014 436137 126082 436193
rect 126138 436137 126208 436193
rect 125888 436069 126208 436137
rect 125888 436013 125958 436069
rect 126014 436013 126082 436069
rect 126138 436013 126208 436069
rect 95168 435889 95238 435945
rect 95294 435889 95362 435945
rect 95418 435889 95488 435945
rect 95168 435826 95488 435889
rect 125888 435945 126208 436013
rect 129154 436378 129774 453922
rect 129154 436322 129250 436378
rect 129306 436322 129374 436378
rect 129430 436322 129498 436378
rect 129554 436322 129622 436378
rect 129678 436322 129774 436378
rect 129154 436254 129774 436322
rect 129154 436198 129250 436254
rect 129306 436198 129374 436254
rect 129430 436198 129498 436254
rect 129554 436198 129622 436254
rect 129678 436198 129774 436254
rect 129154 436130 129774 436198
rect 129154 436074 129250 436130
rect 129306 436074 129374 436130
rect 129430 436074 129498 436130
rect 129554 436074 129622 436130
rect 129678 436074 129774 436130
rect 129154 436006 129774 436074
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 514350 133494 531922
rect 132874 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 133494 514350
rect 132874 514226 133494 514294
rect 132874 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 133494 514226
rect 132874 514102 133494 514170
rect 132874 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 133494 514102
rect 132874 513978 133494 514046
rect 132874 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 133494 513978
rect 132874 496350 133494 513922
rect 132874 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 133494 496350
rect 132874 496226 133494 496294
rect 132874 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 133494 496226
rect 132874 496102 133494 496170
rect 132874 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 133494 496102
rect 132874 495978 133494 496046
rect 132874 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 133494 495978
rect 132874 478350 133494 495922
rect 132874 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 133494 478350
rect 132874 478226 133494 478294
rect 132874 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 133494 478226
rect 132874 478102 133494 478170
rect 132874 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 133494 478102
rect 132874 477978 133494 478046
rect 132874 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 133494 477978
rect 132874 460350 133494 477922
rect 132874 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 133494 460350
rect 132874 460226 133494 460294
rect 132874 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 133494 460226
rect 132874 460102 133494 460170
rect 132874 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 133494 460102
rect 132874 459978 133494 460046
rect 132874 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 133494 459978
rect 132874 442350 133494 459922
rect 132874 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 133494 442350
rect 132874 442226 133494 442294
rect 132874 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 133494 442226
rect 132874 442102 133494 442170
rect 132874 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 133494 442102
rect 132874 441978 133494 442046
rect 132874 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 133494 441978
rect 132874 436006 133494 441922
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 526350 147774 543922
rect 147154 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 147774 526350
rect 147154 526226 147774 526294
rect 147154 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 147774 526226
rect 147154 526102 147774 526170
rect 147154 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 147774 526102
rect 147154 525978 147774 526046
rect 147154 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 147774 525978
rect 147154 508350 147774 525922
rect 147154 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 147774 508350
rect 147154 508226 147774 508294
rect 147154 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 147774 508226
rect 147154 508102 147774 508170
rect 147154 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 147774 508102
rect 147154 507978 147774 508046
rect 147154 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 147774 507978
rect 147154 490350 147774 507922
rect 147154 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 147774 490350
rect 147154 490226 147774 490294
rect 147154 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 147774 490226
rect 147154 490102 147774 490170
rect 147154 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 147774 490102
rect 147154 489978 147774 490046
rect 147154 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 147774 489978
rect 147154 472350 147774 489922
rect 147154 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 147774 472350
rect 147154 472226 147774 472294
rect 147154 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 147774 472226
rect 147154 472102 147774 472170
rect 147154 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 147774 472102
rect 147154 471978 147774 472046
rect 147154 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 147774 471978
rect 147154 454350 147774 471922
rect 147154 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 147774 454350
rect 147154 454226 147774 454294
rect 147154 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 147774 454226
rect 147154 454102 147774 454170
rect 147154 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 147774 454102
rect 147154 453978 147774 454046
rect 147154 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 147774 453978
rect 147154 436378 147774 453922
rect 147154 436322 147250 436378
rect 147306 436322 147374 436378
rect 147430 436322 147498 436378
rect 147554 436322 147622 436378
rect 147678 436322 147774 436378
rect 147154 436254 147774 436322
rect 147154 436198 147250 436254
rect 147306 436198 147374 436254
rect 147430 436198 147498 436254
rect 147554 436198 147622 436254
rect 147678 436198 147774 436254
rect 147154 436130 147774 436198
rect 147154 436074 147250 436130
rect 147306 436074 147374 436130
rect 147430 436074 147498 436130
rect 147554 436074 147622 436130
rect 147678 436074 147774 436130
rect 147154 436006 147774 436074
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 514350 151494 531922
rect 150874 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 151494 514350
rect 150874 514226 151494 514294
rect 150874 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 151494 514226
rect 150874 514102 151494 514170
rect 150874 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 151494 514102
rect 150874 513978 151494 514046
rect 150874 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 151494 513978
rect 150874 496350 151494 513922
rect 150874 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 151494 496350
rect 150874 496226 151494 496294
rect 150874 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 151494 496226
rect 150874 496102 151494 496170
rect 150874 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 151494 496102
rect 150874 495978 151494 496046
rect 150874 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 151494 495978
rect 150874 478350 151494 495922
rect 150874 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 151494 478350
rect 150874 478226 151494 478294
rect 150874 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 151494 478226
rect 150874 478102 151494 478170
rect 150874 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 151494 478102
rect 150874 477978 151494 478046
rect 150874 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 151494 477978
rect 150874 460350 151494 477922
rect 150874 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 151494 460350
rect 150874 460226 151494 460294
rect 150874 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 151494 460226
rect 150874 460102 151494 460170
rect 150874 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 151494 460102
rect 150874 459978 151494 460046
rect 150874 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 151494 459978
rect 150874 442350 151494 459922
rect 150874 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 151494 442350
rect 150874 442226 151494 442294
rect 150874 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 151494 442226
rect 150874 442102 151494 442170
rect 150874 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 151494 442102
rect 150874 441978 151494 442046
rect 150874 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 151494 441978
rect 150874 436006 151494 441922
rect 165154 597212 165774 598268
rect 165154 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 165774 597212
rect 165154 597088 165774 597156
rect 165154 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 165774 597088
rect 165154 596964 165774 597032
rect 165154 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 165774 596964
rect 165154 596840 165774 596908
rect 165154 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 165774 596840
rect 165154 580350 165774 596784
rect 165154 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 165774 580350
rect 165154 580226 165774 580294
rect 165154 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 165774 580226
rect 165154 580102 165774 580170
rect 165154 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 165774 580102
rect 165154 579978 165774 580046
rect 165154 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 165774 579978
rect 165154 562350 165774 579922
rect 165154 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 165774 562350
rect 165154 562226 165774 562294
rect 165154 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 165774 562226
rect 165154 562102 165774 562170
rect 165154 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 165774 562102
rect 165154 561978 165774 562046
rect 165154 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 165774 561978
rect 165154 544350 165774 561922
rect 165154 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 165774 544350
rect 165154 544226 165774 544294
rect 165154 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 165774 544226
rect 165154 544102 165774 544170
rect 165154 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 165774 544102
rect 165154 543978 165774 544046
rect 165154 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 165774 543978
rect 165154 526350 165774 543922
rect 165154 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 165774 526350
rect 165154 526226 165774 526294
rect 165154 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 165774 526226
rect 165154 526102 165774 526170
rect 165154 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 165774 526102
rect 165154 525978 165774 526046
rect 165154 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 165774 525978
rect 165154 508350 165774 525922
rect 165154 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 165774 508350
rect 165154 508226 165774 508294
rect 165154 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 165774 508226
rect 165154 508102 165774 508170
rect 165154 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 165774 508102
rect 165154 507978 165774 508046
rect 165154 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 165774 507978
rect 165154 490350 165774 507922
rect 165154 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 165774 490350
rect 165154 490226 165774 490294
rect 165154 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 165774 490226
rect 165154 490102 165774 490170
rect 165154 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 165774 490102
rect 165154 489978 165774 490046
rect 165154 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 165774 489978
rect 165154 472350 165774 489922
rect 165154 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 165774 472350
rect 165154 472226 165774 472294
rect 165154 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 165774 472226
rect 165154 472102 165774 472170
rect 165154 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 165774 472102
rect 165154 471978 165774 472046
rect 165154 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 165774 471978
rect 165154 454350 165774 471922
rect 165154 454294 165250 454350
rect 165306 454294 165374 454350
rect 165430 454294 165498 454350
rect 165554 454294 165622 454350
rect 165678 454294 165774 454350
rect 165154 454226 165774 454294
rect 165154 454170 165250 454226
rect 165306 454170 165374 454226
rect 165430 454170 165498 454226
rect 165554 454170 165622 454226
rect 165678 454170 165774 454226
rect 165154 454102 165774 454170
rect 165154 454046 165250 454102
rect 165306 454046 165374 454102
rect 165430 454046 165498 454102
rect 165554 454046 165622 454102
rect 165678 454046 165774 454102
rect 165154 453978 165774 454046
rect 165154 453922 165250 453978
rect 165306 453922 165374 453978
rect 165430 453922 165498 453978
rect 165554 453922 165622 453978
rect 165678 453922 165774 453978
rect 156608 436317 156928 436380
rect 156608 436261 156678 436317
rect 156734 436261 156802 436317
rect 156858 436261 156928 436317
rect 156608 436193 156928 436261
rect 156608 436137 156678 436193
rect 156734 436137 156802 436193
rect 156858 436137 156928 436193
rect 156608 436069 156928 436137
rect 156608 436013 156678 436069
rect 156734 436013 156802 436069
rect 156858 436013 156928 436069
rect 125888 435889 125958 435945
rect 126014 435889 126082 435945
rect 126138 435889 126208 435945
rect 125888 435826 126208 435889
rect 156608 435945 156928 436013
rect 165154 436378 165774 453922
rect 165154 436322 165250 436378
rect 165306 436322 165374 436378
rect 165430 436322 165498 436378
rect 165554 436322 165622 436378
rect 165678 436322 165774 436378
rect 165154 436254 165774 436322
rect 165154 436198 165250 436254
rect 165306 436198 165374 436254
rect 165430 436198 165498 436254
rect 165554 436198 165622 436254
rect 165678 436198 165774 436254
rect 165154 436130 165774 436198
rect 165154 436074 165250 436130
rect 165306 436074 165374 436130
rect 165430 436074 165498 436130
rect 165554 436074 165622 436130
rect 165678 436074 165774 436130
rect 165154 436006 165774 436074
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 514350 169494 531922
rect 168874 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 169494 514350
rect 168874 514226 169494 514294
rect 168874 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 169494 514226
rect 168874 514102 169494 514170
rect 168874 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 169494 514102
rect 168874 513978 169494 514046
rect 168874 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 169494 513978
rect 168874 496350 169494 513922
rect 168874 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 169494 496350
rect 168874 496226 169494 496294
rect 168874 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 169494 496226
rect 168874 496102 169494 496170
rect 168874 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 169494 496102
rect 168874 495978 169494 496046
rect 168874 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 169494 495978
rect 168874 478350 169494 495922
rect 168874 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 169494 478350
rect 168874 478226 169494 478294
rect 168874 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 169494 478226
rect 168874 478102 169494 478170
rect 168874 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 169494 478102
rect 168874 477978 169494 478046
rect 168874 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 169494 477978
rect 168874 460350 169494 477922
rect 168874 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 169494 460350
rect 168874 460226 169494 460294
rect 168874 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 169494 460226
rect 168874 460102 169494 460170
rect 168874 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 169494 460102
rect 168874 459978 169494 460046
rect 168874 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 169494 459978
rect 168874 442350 169494 459922
rect 168874 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 169494 442350
rect 168874 442226 169494 442294
rect 168874 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 169494 442226
rect 168874 442102 169494 442170
rect 168874 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 169494 442102
rect 168874 441978 169494 442046
rect 168874 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 169494 441978
rect 168874 436006 169494 441922
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 526350 183774 543922
rect 183154 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 183774 526350
rect 183154 526226 183774 526294
rect 183154 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 183774 526226
rect 183154 526102 183774 526170
rect 183154 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 183774 526102
rect 183154 525978 183774 526046
rect 183154 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 183774 525978
rect 183154 508350 183774 525922
rect 183154 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 183774 508350
rect 183154 508226 183774 508294
rect 183154 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 183774 508226
rect 183154 508102 183774 508170
rect 183154 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 183774 508102
rect 183154 507978 183774 508046
rect 183154 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 183774 507978
rect 183154 490350 183774 507922
rect 183154 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 183774 490350
rect 183154 490226 183774 490294
rect 183154 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 183774 490226
rect 183154 490102 183774 490170
rect 183154 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 183774 490102
rect 183154 489978 183774 490046
rect 183154 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 183774 489978
rect 183154 472350 183774 489922
rect 183154 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 183774 472350
rect 183154 472226 183774 472294
rect 183154 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 183774 472226
rect 183154 472102 183774 472170
rect 183154 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 183774 472102
rect 183154 471978 183774 472046
rect 183154 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 183774 471978
rect 183154 454350 183774 471922
rect 183154 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 183774 454350
rect 183154 454226 183774 454294
rect 183154 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 183774 454226
rect 183154 454102 183774 454170
rect 183154 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 183774 454102
rect 183154 453978 183774 454046
rect 183154 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 183774 453978
rect 183154 436378 183774 453922
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 514350 187494 531922
rect 186874 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 187494 514350
rect 186874 514226 187494 514294
rect 186874 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 187494 514226
rect 186874 514102 187494 514170
rect 186874 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 187494 514102
rect 186874 513978 187494 514046
rect 186874 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 187494 513978
rect 186874 496350 187494 513922
rect 186874 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 187494 496350
rect 186874 496226 187494 496294
rect 186874 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 187494 496226
rect 186874 496102 187494 496170
rect 186874 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 187494 496102
rect 186874 495978 187494 496046
rect 186874 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 187494 495978
rect 186874 478350 187494 495922
rect 186874 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 187494 478350
rect 186874 478226 187494 478294
rect 186874 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 187494 478226
rect 186874 478102 187494 478170
rect 186874 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 187494 478102
rect 186874 477978 187494 478046
rect 186874 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 187494 477978
rect 186874 460350 187494 477922
rect 186874 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 187494 460350
rect 186874 460226 187494 460294
rect 186874 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 187494 460226
rect 186874 460102 187494 460170
rect 186874 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 187494 460102
rect 186874 459978 187494 460046
rect 186874 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 187494 459978
rect 186874 442350 187494 459922
rect 186874 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 187494 442350
rect 186874 442226 187494 442294
rect 186874 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 187494 442226
rect 186874 442102 187494 442170
rect 186874 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 187494 442102
rect 186874 441978 187494 442046
rect 186874 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 187494 441978
rect 186874 438436 187494 441922
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 526350 201774 543922
rect 201154 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 201774 526350
rect 201154 526226 201774 526294
rect 201154 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 201774 526226
rect 201154 526102 201774 526170
rect 201154 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 201774 526102
rect 201154 525978 201774 526046
rect 201154 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 201774 525978
rect 201154 508350 201774 525922
rect 201154 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 201774 508350
rect 201154 508226 201774 508294
rect 201154 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 201774 508226
rect 201154 508102 201774 508170
rect 201154 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 201774 508102
rect 201154 507978 201774 508046
rect 201154 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 201774 507978
rect 201154 490350 201774 507922
rect 201154 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 201774 490350
rect 201154 490226 201774 490294
rect 201154 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 201774 490226
rect 201154 490102 201774 490170
rect 201154 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 201774 490102
rect 201154 489978 201774 490046
rect 201154 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 201774 489978
rect 201154 472350 201774 489922
rect 201154 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 201774 472350
rect 201154 472226 201774 472294
rect 201154 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 201774 472226
rect 201154 472102 201774 472170
rect 201154 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 201774 472102
rect 201154 471978 201774 472046
rect 201154 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 201774 471978
rect 201154 454350 201774 471922
rect 201154 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 201774 454350
rect 201154 454226 201774 454294
rect 201154 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 201774 454226
rect 201154 454102 201774 454170
rect 201154 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 201774 454102
rect 201154 453978 201774 454046
rect 201154 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 201774 453978
rect 183154 436322 183250 436378
rect 183306 436322 183374 436378
rect 183430 436322 183498 436378
rect 183554 436322 183622 436378
rect 183678 436322 183774 436378
rect 183154 436254 183774 436322
rect 183154 436198 183250 436254
rect 183306 436198 183374 436254
rect 183430 436198 183498 436254
rect 183554 436198 183622 436254
rect 183678 436198 183774 436254
rect 183154 436130 183774 436198
rect 183154 436074 183250 436130
rect 183306 436074 183374 436130
rect 183430 436074 183498 436130
rect 183554 436074 183622 436130
rect 183678 436074 183774 436130
rect 183154 436006 183774 436074
rect 187328 436317 187648 436380
rect 187328 436261 187398 436317
rect 187454 436261 187522 436317
rect 187578 436261 187648 436317
rect 187328 436193 187648 436261
rect 187328 436137 187398 436193
rect 187454 436137 187522 436193
rect 187578 436137 187648 436193
rect 187328 436069 187648 436137
rect 187328 436013 187398 436069
rect 187454 436013 187522 436069
rect 187578 436013 187648 436069
rect 156608 435889 156678 435945
rect 156734 435889 156802 435945
rect 156858 435889 156928 435945
rect 156608 435826 156928 435889
rect 187328 435945 187648 436013
rect 201154 436378 201774 453922
rect 201154 436322 201250 436378
rect 201306 436322 201374 436378
rect 201430 436322 201498 436378
rect 201554 436322 201622 436378
rect 201678 436322 201774 436378
rect 201154 436254 201774 436322
rect 201154 436198 201250 436254
rect 201306 436198 201374 436254
rect 201430 436198 201498 436254
rect 201554 436198 201622 436254
rect 201678 436198 201774 436254
rect 201154 436130 201774 436198
rect 201154 436074 201250 436130
rect 201306 436074 201374 436130
rect 201430 436074 201498 436130
rect 201554 436074 201622 436130
rect 201678 436074 201774 436130
rect 201154 436006 201774 436074
rect 204874 598172 205494 598268
rect 204874 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 205494 598172
rect 204874 598048 205494 598116
rect 204874 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 205494 598048
rect 204874 597924 205494 597992
rect 204874 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 205494 597924
rect 204874 597800 205494 597868
rect 204874 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 205494 597800
rect 204874 586350 205494 597744
rect 204874 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 205494 586350
rect 204874 586226 205494 586294
rect 204874 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 205494 586226
rect 204874 586102 205494 586170
rect 204874 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 205494 586102
rect 204874 585978 205494 586046
rect 204874 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 205494 585978
rect 204874 568350 205494 585922
rect 204874 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 205494 568350
rect 204874 568226 205494 568294
rect 204874 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 205494 568226
rect 204874 568102 205494 568170
rect 204874 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 205494 568102
rect 204874 567978 205494 568046
rect 204874 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 205494 567978
rect 204874 550350 205494 567922
rect 204874 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 205494 550350
rect 204874 550226 205494 550294
rect 204874 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 205494 550226
rect 204874 550102 205494 550170
rect 204874 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 205494 550102
rect 204874 549978 205494 550046
rect 204874 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 205494 549978
rect 204874 532350 205494 549922
rect 204874 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 205494 532350
rect 204874 532226 205494 532294
rect 204874 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 205494 532226
rect 204874 532102 205494 532170
rect 204874 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 205494 532102
rect 204874 531978 205494 532046
rect 204874 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 205494 531978
rect 204874 514350 205494 531922
rect 204874 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 205494 514350
rect 204874 514226 205494 514294
rect 204874 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 205494 514226
rect 204874 514102 205494 514170
rect 204874 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 205494 514102
rect 204874 513978 205494 514046
rect 204874 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 205494 513978
rect 204874 496350 205494 513922
rect 204874 496294 204970 496350
rect 205026 496294 205094 496350
rect 205150 496294 205218 496350
rect 205274 496294 205342 496350
rect 205398 496294 205494 496350
rect 204874 496226 205494 496294
rect 204874 496170 204970 496226
rect 205026 496170 205094 496226
rect 205150 496170 205218 496226
rect 205274 496170 205342 496226
rect 205398 496170 205494 496226
rect 204874 496102 205494 496170
rect 204874 496046 204970 496102
rect 205026 496046 205094 496102
rect 205150 496046 205218 496102
rect 205274 496046 205342 496102
rect 205398 496046 205494 496102
rect 204874 495978 205494 496046
rect 204874 495922 204970 495978
rect 205026 495922 205094 495978
rect 205150 495922 205218 495978
rect 205274 495922 205342 495978
rect 205398 495922 205494 495978
rect 204874 478350 205494 495922
rect 204874 478294 204970 478350
rect 205026 478294 205094 478350
rect 205150 478294 205218 478350
rect 205274 478294 205342 478350
rect 205398 478294 205494 478350
rect 204874 478226 205494 478294
rect 204874 478170 204970 478226
rect 205026 478170 205094 478226
rect 205150 478170 205218 478226
rect 205274 478170 205342 478226
rect 205398 478170 205494 478226
rect 204874 478102 205494 478170
rect 204874 478046 204970 478102
rect 205026 478046 205094 478102
rect 205150 478046 205218 478102
rect 205274 478046 205342 478102
rect 205398 478046 205494 478102
rect 204874 477978 205494 478046
rect 204874 477922 204970 477978
rect 205026 477922 205094 477978
rect 205150 477922 205218 477978
rect 205274 477922 205342 477978
rect 205398 477922 205494 477978
rect 204874 460350 205494 477922
rect 204874 460294 204970 460350
rect 205026 460294 205094 460350
rect 205150 460294 205218 460350
rect 205274 460294 205342 460350
rect 205398 460294 205494 460350
rect 204874 460226 205494 460294
rect 204874 460170 204970 460226
rect 205026 460170 205094 460226
rect 205150 460170 205218 460226
rect 205274 460170 205342 460226
rect 205398 460170 205494 460226
rect 204874 460102 205494 460170
rect 204874 460046 204970 460102
rect 205026 460046 205094 460102
rect 205150 460046 205218 460102
rect 205274 460046 205342 460102
rect 205398 460046 205494 460102
rect 204874 459978 205494 460046
rect 204874 459922 204970 459978
rect 205026 459922 205094 459978
rect 205150 459922 205218 459978
rect 205274 459922 205342 459978
rect 205398 459922 205494 459978
rect 204874 442350 205494 459922
rect 204874 442294 204970 442350
rect 205026 442294 205094 442350
rect 205150 442294 205218 442350
rect 205274 442294 205342 442350
rect 205398 442294 205494 442350
rect 204874 442226 205494 442294
rect 204874 442170 204970 442226
rect 205026 442170 205094 442226
rect 205150 442170 205218 442226
rect 205274 442170 205342 442226
rect 205398 442170 205494 442226
rect 204874 442102 205494 442170
rect 204874 442046 204970 442102
rect 205026 442046 205094 442102
rect 205150 442046 205218 442102
rect 205274 442046 205342 442102
rect 205398 442046 205494 442102
rect 204874 441978 205494 442046
rect 204874 441922 204970 441978
rect 205026 441922 205094 441978
rect 205150 441922 205218 441978
rect 205274 441922 205342 441978
rect 205398 441922 205494 441978
rect 204874 436006 205494 441922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 526350 219774 543922
rect 219154 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 219774 526350
rect 219154 526226 219774 526294
rect 219154 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 219774 526226
rect 219154 526102 219774 526170
rect 219154 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 219774 526102
rect 219154 525978 219774 526046
rect 219154 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 219774 525978
rect 219154 508350 219774 525922
rect 219154 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 219774 508350
rect 219154 508226 219774 508294
rect 219154 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 219774 508226
rect 219154 508102 219774 508170
rect 219154 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 219774 508102
rect 219154 507978 219774 508046
rect 219154 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 219774 507978
rect 219154 490350 219774 507922
rect 219154 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 219774 490350
rect 219154 490226 219774 490294
rect 219154 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 219774 490226
rect 219154 490102 219774 490170
rect 219154 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 219774 490102
rect 219154 489978 219774 490046
rect 219154 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 219774 489978
rect 219154 472350 219774 489922
rect 219154 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 219774 472350
rect 219154 472226 219774 472294
rect 219154 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 219774 472226
rect 219154 472102 219774 472170
rect 219154 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 219774 472102
rect 219154 471978 219774 472046
rect 219154 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 219774 471978
rect 219154 454350 219774 471922
rect 219154 454294 219250 454350
rect 219306 454294 219374 454350
rect 219430 454294 219498 454350
rect 219554 454294 219622 454350
rect 219678 454294 219774 454350
rect 219154 454226 219774 454294
rect 219154 454170 219250 454226
rect 219306 454170 219374 454226
rect 219430 454170 219498 454226
rect 219554 454170 219622 454226
rect 219678 454170 219774 454226
rect 219154 454102 219774 454170
rect 219154 454046 219250 454102
rect 219306 454046 219374 454102
rect 219430 454046 219498 454102
rect 219554 454046 219622 454102
rect 219678 454046 219774 454102
rect 219154 453978 219774 454046
rect 219154 453922 219250 453978
rect 219306 453922 219374 453978
rect 219430 453922 219498 453978
rect 219554 453922 219622 453978
rect 219678 453922 219774 453978
rect 218048 436317 218368 436380
rect 218048 436261 218118 436317
rect 218174 436261 218242 436317
rect 218298 436261 218368 436317
rect 218048 436193 218368 436261
rect 218048 436137 218118 436193
rect 218174 436137 218242 436193
rect 218298 436137 218368 436193
rect 218048 436069 218368 436137
rect 218048 436013 218118 436069
rect 218174 436013 218242 436069
rect 218298 436013 218368 436069
rect 187328 435889 187398 435945
rect 187454 435889 187522 435945
rect 187578 435889 187648 435945
rect 187328 435826 187648 435889
rect 218048 435945 218368 436013
rect 219154 436378 219774 453922
rect 219154 436322 219250 436378
rect 219306 436322 219374 436378
rect 219430 436322 219498 436378
rect 219554 436322 219622 436378
rect 219678 436322 219774 436378
rect 219154 436254 219774 436322
rect 219154 436198 219250 436254
rect 219306 436198 219374 436254
rect 219430 436198 219498 436254
rect 219554 436198 219622 436254
rect 219678 436198 219774 436254
rect 219154 436130 219774 436198
rect 219154 436074 219250 436130
rect 219306 436074 219374 436130
rect 219430 436074 219498 436130
rect 219554 436074 219622 436130
rect 219678 436074 219774 436130
rect 219154 436006 219774 436074
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 514350 223494 531922
rect 222874 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 223494 514350
rect 222874 514226 223494 514294
rect 222874 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 223494 514226
rect 222874 514102 223494 514170
rect 222874 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 223494 514102
rect 222874 513978 223494 514046
rect 222874 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 223494 513978
rect 222874 496350 223494 513922
rect 222874 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 223494 496350
rect 222874 496226 223494 496294
rect 222874 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 223494 496226
rect 222874 496102 223494 496170
rect 222874 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 223494 496102
rect 222874 495978 223494 496046
rect 222874 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 223494 495978
rect 222874 478350 223494 495922
rect 222874 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 223494 478350
rect 222874 478226 223494 478294
rect 222874 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 223494 478226
rect 222874 478102 223494 478170
rect 222874 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 223494 478102
rect 222874 477978 223494 478046
rect 222874 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 223494 477978
rect 222874 460350 223494 477922
rect 222874 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 223494 460350
rect 222874 460226 223494 460294
rect 222874 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 223494 460226
rect 222874 460102 223494 460170
rect 222874 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 223494 460102
rect 222874 459978 223494 460046
rect 222874 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 223494 459978
rect 222874 442350 223494 459922
rect 222874 442294 222970 442350
rect 223026 442294 223094 442350
rect 223150 442294 223218 442350
rect 223274 442294 223342 442350
rect 223398 442294 223494 442350
rect 222874 442226 223494 442294
rect 222874 442170 222970 442226
rect 223026 442170 223094 442226
rect 223150 442170 223218 442226
rect 223274 442170 223342 442226
rect 223398 442170 223494 442226
rect 222874 442102 223494 442170
rect 222874 442046 222970 442102
rect 223026 442046 223094 442102
rect 223150 442046 223218 442102
rect 223274 442046 223342 442102
rect 223398 442046 223494 442102
rect 222874 441978 223494 442046
rect 222874 441922 222970 441978
rect 223026 441922 223094 441978
rect 223150 441922 223218 441978
rect 223274 441922 223342 441978
rect 223398 441922 223494 441978
rect 222874 436006 223494 441922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 526350 237774 543922
rect 237154 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 237774 526350
rect 237154 526226 237774 526294
rect 237154 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 237774 526226
rect 237154 526102 237774 526170
rect 237154 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 237774 526102
rect 237154 525978 237774 526046
rect 237154 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 237774 525978
rect 237154 508350 237774 525922
rect 237154 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 237774 508350
rect 237154 508226 237774 508294
rect 237154 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 237774 508226
rect 237154 508102 237774 508170
rect 237154 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 237774 508102
rect 237154 507978 237774 508046
rect 237154 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 237774 507978
rect 237154 490350 237774 507922
rect 237154 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 237774 490350
rect 237154 490226 237774 490294
rect 237154 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 237774 490226
rect 237154 490102 237774 490170
rect 237154 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 237774 490102
rect 237154 489978 237774 490046
rect 237154 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 237774 489978
rect 237154 472350 237774 489922
rect 237154 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 237774 472350
rect 237154 472226 237774 472294
rect 237154 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 237774 472226
rect 237154 472102 237774 472170
rect 237154 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 237774 472102
rect 237154 471978 237774 472046
rect 237154 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 237774 471978
rect 237154 454350 237774 471922
rect 237154 454294 237250 454350
rect 237306 454294 237374 454350
rect 237430 454294 237498 454350
rect 237554 454294 237622 454350
rect 237678 454294 237774 454350
rect 237154 454226 237774 454294
rect 237154 454170 237250 454226
rect 237306 454170 237374 454226
rect 237430 454170 237498 454226
rect 237554 454170 237622 454226
rect 237678 454170 237774 454226
rect 237154 454102 237774 454170
rect 237154 454046 237250 454102
rect 237306 454046 237374 454102
rect 237430 454046 237498 454102
rect 237554 454046 237622 454102
rect 237678 454046 237774 454102
rect 237154 453978 237774 454046
rect 237154 453922 237250 453978
rect 237306 453922 237374 453978
rect 237430 453922 237498 453978
rect 237554 453922 237622 453978
rect 237678 453922 237774 453978
rect 237154 436378 237774 453922
rect 237154 436322 237250 436378
rect 237306 436322 237374 436378
rect 237430 436322 237498 436378
rect 237554 436322 237622 436378
rect 237678 436322 237774 436378
rect 237154 436254 237774 436322
rect 237154 436198 237250 436254
rect 237306 436198 237374 436254
rect 237430 436198 237498 436254
rect 237554 436198 237622 436254
rect 237678 436198 237774 436254
rect 237154 436130 237774 436198
rect 237154 436074 237250 436130
rect 237306 436074 237374 436130
rect 237430 436074 237498 436130
rect 237554 436074 237622 436130
rect 237678 436074 237774 436130
rect 237154 436006 237774 436074
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 514350 241494 531922
rect 240874 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 241494 514350
rect 240874 514226 241494 514294
rect 240874 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 241494 514226
rect 240874 514102 241494 514170
rect 240874 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 241494 514102
rect 240874 513978 241494 514046
rect 240874 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 241494 513978
rect 240874 496350 241494 513922
rect 240874 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 241494 496350
rect 240874 496226 241494 496294
rect 240874 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 241494 496226
rect 240874 496102 241494 496170
rect 240874 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 241494 496102
rect 240874 495978 241494 496046
rect 240874 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 241494 495978
rect 240874 478350 241494 495922
rect 240874 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 241494 478350
rect 240874 478226 241494 478294
rect 240874 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 241494 478226
rect 240874 478102 241494 478170
rect 240874 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 241494 478102
rect 240874 477978 241494 478046
rect 240874 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 241494 477978
rect 240874 460350 241494 477922
rect 240874 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 241494 460350
rect 240874 460226 241494 460294
rect 240874 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 241494 460226
rect 240874 460102 241494 460170
rect 240874 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 241494 460102
rect 240874 459978 241494 460046
rect 240874 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 241494 459978
rect 240874 442350 241494 459922
rect 240874 442294 240970 442350
rect 241026 442294 241094 442350
rect 241150 442294 241218 442350
rect 241274 442294 241342 442350
rect 241398 442294 241494 442350
rect 240874 442226 241494 442294
rect 240874 442170 240970 442226
rect 241026 442170 241094 442226
rect 241150 442170 241218 442226
rect 241274 442170 241342 442226
rect 241398 442170 241494 442226
rect 240874 442102 241494 442170
rect 240874 442046 240970 442102
rect 241026 442046 241094 442102
rect 241150 442046 241218 442102
rect 241274 442046 241342 442102
rect 241398 442046 241494 442102
rect 240874 441978 241494 442046
rect 240874 441922 240970 441978
rect 241026 441922 241094 441978
rect 241150 441922 241218 441978
rect 241274 441922 241342 441978
rect 241398 441922 241494 441978
rect 240874 436006 241494 441922
rect 255154 597212 255774 598268
rect 255154 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 255774 597212
rect 255154 597088 255774 597156
rect 255154 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 255774 597088
rect 255154 596964 255774 597032
rect 255154 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 255774 596964
rect 255154 596840 255774 596908
rect 255154 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 255774 596840
rect 255154 580350 255774 596784
rect 255154 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 255774 580350
rect 255154 580226 255774 580294
rect 255154 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 255774 580226
rect 255154 580102 255774 580170
rect 255154 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 255774 580102
rect 255154 579978 255774 580046
rect 255154 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 255774 579978
rect 255154 562350 255774 579922
rect 255154 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 255774 562350
rect 255154 562226 255774 562294
rect 255154 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 255774 562226
rect 255154 562102 255774 562170
rect 255154 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 255774 562102
rect 255154 561978 255774 562046
rect 255154 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 255774 561978
rect 255154 544350 255774 561922
rect 255154 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 255774 544350
rect 255154 544226 255774 544294
rect 255154 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 255774 544226
rect 255154 544102 255774 544170
rect 255154 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 255774 544102
rect 255154 543978 255774 544046
rect 255154 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 255774 543978
rect 255154 526350 255774 543922
rect 255154 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 255774 526350
rect 255154 526226 255774 526294
rect 255154 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 255774 526226
rect 255154 526102 255774 526170
rect 255154 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 255774 526102
rect 255154 525978 255774 526046
rect 255154 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 255774 525978
rect 255154 508350 255774 525922
rect 255154 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 255774 508350
rect 255154 508226 255774 508294
rect 255154 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 255774 508226
rect 255154 508102 255774 508170
rect 255154 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 255774 508102
rect 255154 507978 255774 508046
rect 255154 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 255774 507978
rect 255154 490350 255774 507922
rect 255154 490294 255250 490350
rect 255306 490294 255374 490350
rect 255430 490294 255498 490350
rect 255554 490294 255622 490350
rect 255678 490294 255774 490350
rect 255154 490226 255774 490294
rect 255154 490170 255250 490226
rect 255306 490170 255374 490226
rect 255430 490170 255498 490226
rect 255554 490170 255622 490226
rect 255678 490170 255774 490226
rect 255154 490102 255774 490170
rect 255154 490046 255250 490102
rect 255306 490046 255374 490102
rect 255430 490046 255498 490102
rect 255554 490046 255622 490102
rect 255678 490046 255774 490102
rect 255154 489978 255774 490046
rect 255154 489922 255250 489978
rect 255306 489922 255374 489978
rect 255430 489922 255498 489978
rect 255554 489922 255622 489978
rect 255678 489922 255774 489978
rect 255154 472350 255774 489922
rect 255154 472294 255250 472350
rect 255306 472294 255374 472350
rect 255430 472294 255498 472350
rect 255554 472294 255622 472350
rect 255678 472294 255774 472350
rect 255154 472226 255774 472294
rect 255154 472170 255250 472226
rect 255306 472170 255374 472226
rect 255430 472170 255498 472226
rect 255554 472170 255622 472226
rect 255678 472170 255774 472226
rect 255154 472102 255774 472170
rect 255154 472046 255250 472102
rect 255306 472046 255374 472102
rect 255430 472046 255498 472102
rect 255554 472046 255622 472102
rect 255678 472046 255774 472102
rect 255154 471978 255774 472046
rect 255154 471922 255250 471978
rect 255306 471922 255374 471978
rect 255430 471922 255498 471978
rect 255554 471922 255622 471978
rect 255678 471922 255774 471978
rect 255154 454350 255774 471922
rect 255154 454294 255250 454350
rect 255306 454294 255374 454350
rect 255430 454294 255498 454350
rect 255554 454294 255622 454350
rect 255678 454294 255774 454350
rect 255154 454226 255774 454294
rect 255154 454170 255250 454226
rect 255306 454170 255374 454226
rect 255430 454170 255498 454226
rect 255554 454170 255622 454226
rect 255678 454170 255774 454226
rect 255154 454102 255774 454170
rect 255154 454046 255250 454102
rect 255306 454046 255374 454102
rect 255430 454046 255498 454102
rect 255554 454046 255622 454102
rect 255678 454046 255774 454102
rect 255154 453978 255774 454046
rect 255154 453922 255250 453978
rect 255306 453922 255374 453978
rect 255430 453922 255498 453978
rect 255554 453922 255622 453978
rect 255678 453922 255774 453978
rect 248768 436317 249088 436380
rect 248768 436261 248838 436317
rect 248894 436261 248962 436317
rect 249018 436261 249088 436317
rect 248768 436193 249088 436261
rect 248768 436137 248838 436193
rect 248894 436137 248962 436193
rect 249018 436137 249088 436193
rect 248768 436069 249088 436137
rect 248768 436013 248838 436069
rect 248894 436013 248962 436069
rect 249018 436013 249088 436069
rect 218048 435889 218118 435945
rect 218174 435889 218242 435945
rect 218298 435889 218368 435945
rect 218048 435826 218368 435889
rect 248768 435945 249088 436013
rect 255154 436378 255774 453922
rect 255154 436322 255250 436378
rect 255306 436322 255374 436378
rect 255430 436322 255498 436378
rect 255554 436322 255622 436378
rect 255678 436322 255774 436378
rect 255154 436254 255774 436322
rect 255154 436198 255250 436254
rect 255306 436198 255374 436254
rect 255430 436198 255498 436254
rect 255554 436198 255622 436254
rect 255678 436198 255774 436254
rect 255154 436130 255774 436198
rect 255154 436074 255250 436130
rect 255306 436074 255374 436130
rect 255430 436074 255498 436130
rect 255554 436074 255622 436130
rect 255678 436074 255774 436130
rect 255154 436006 255774 436074
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 514350 259494 531922
rect 258874 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 259494 514350
rect 258874 514226 259494 514294
rect 258874 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 259494 514226
rect 258874 514102 259494 514170
rect 258874 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 259494 514102
rect 258874 513978 259494 514046
rect 258874 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 259494 513978
rect 258874 496350 259494 513922
rect 258874 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 259494 496350
rect 258874 496226 259494 496294
rect 258874 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 259494 496226
rect 258874 496102 259494 496170
rect 258874 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 259494 496102
rect 258874 495978 259494 496046
rect 258874 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 259494 495978
rect 258874 478350 259494 495922
rect 258874 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 259494 478350
rect 258874 478226 259494 478294
rect 258874 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 259494 478226
rect 258874 478102 259494 478170
rect 258874 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 259494 478102
rect 258874 477978 259494 478046
rect 258874 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 259494 477978
rect 258874 460350 259494 477922
rect 258874 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 259494 460350
rect 258874 460226 259494 460294
rect 258874 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 259494 460226
rect 258874 460102 259494 460170
rect 258874 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 259494 460102
rect 258874 459978 259494 460046
rect 258874 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 259494 459978
rect 258874 442350 259494 459922
rect 258874 442294 258970 442350
rect 259026 442294 259094 442350
rect 259150 442294 259218 442350
rect 259274 442294 259342 442350
rect 259398 442294 259494 442350
rect 258874 442226 259494 442294
rect 258874 442170 258970 442226
rect 259026 442170 259094 442226
rect 259150 442170 259218 442226
rect 259274 442170 259342 442226
rect 259398 442170 259494 442226
rect 258874 442102 259494 442170
rect 258874 442046 258970 442102
rect 259026 442046 259094 442102
rect 259150 442046 259218 442102
rect 259274 442046 259342 442102
rect 259398 442046 259494 442102
rect 258874 441978 259494 442046
rect 258874 441922 258970 441978
rect 259026 441922 259094 441978
rect 259150 441922 259218 441978
rect 259274 441922 259342 441978
rect 259398 441922 259494 441978
rect 258874 436006 259494 441922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 526350 273774 543922
rect 273154 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 273774 526350
rect 273154 526226 273774 526294
rect 273154 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 273774 526226
rect 273154 526102 273774 526170
rect 273154 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 273774 526102
rect 273154 525978 273774 526046
rect 273154 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 273774 525978
rect 273154 508350 273774 525922
rect 273154 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 273774 508350
rect 273154 508226 273774 508294
rect 273154 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 273774 508226
rect 273154 508102 273774 508170
rect 273154 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 273774 508102
rect 273154 507978 273774 508046
rect 273154 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 273774 507978
rect 273154 490350 273774 507922
rect 273154 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 273774 490350
rect 273154 490226 273774 490294
rect 273154 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 273774 490226
rect 273154 490102 273774 490170
rect 273154 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 273774 490102
rect 273154 489978 273774 490046
rect 273154 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 273774 489978
rect 273154 472350 273774 489922
rect 273154 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 273774 472350
rect 273154 472226 273774 472294
rect 273154 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 273774 472226
rect 273154 472102 273774 472170
rect 273154 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 273774 472102
rect 273154 471978 273774 472046
rect 273154 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 273774 471978
rect 273154 454350 273774 471922
rect 273154 454294 273250 454350
rect 273306 454294 273374 454350
rect 273430 454294 273498 454350
rect 273554 454294 273622 454350
rect 273678 454294 273774 454350
rect 273154 454226 273774 454294
rect 273154 454170 273250 454226
rect 273306 454170 273374 454226
rect 273430 454170 273498 454226
rect 273554 454170 273622 454226
rect 273678 454170 273774 454226
rect 273154 454102 273774 454170
rect 273154 454046 273250 454102
rect 273306 454046 273374 454102
rect 273430 454046 273498 454102
rect 273554 454046 273622 454102
rect 273678 454046 273774 454102
rect 273154 453978 273774 454046
rect 273154 453922 273250 453978
rect 273306 453922 273374 453978
rect 273430 453922 273498 453978
rect 273554 453922 273622 453978
rect 273678 453922 273774 453978
rect 273154 436378 273774 453922
rect 273154 436322 273250 436378
rect 273306 436322 273374 436378
rect 273430 436322 273498 436378
rect 273554 436322 273622 436378
rect 273678 436322 273774 436378
rect 273154 436254 273774 436322
rect 273154 436198 273250 436254
rect 273306 436198 273374 436254
rect 273430 436198 273498 436254
rect 273554 436198 273622 436254
rect 273678 436198 273774 436254
rect 273154 436130 273774 436198
rect 273154 436074 273250 436130
rect 273306 436074 273374 436130
rect 273430 436074 273498 436130
rect 273554 436074 273622 436130
rect 273678 436074 273774 436130
rect 273154 436006 273774 436074
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 514350 277494 531922
rect 276874 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 277494 514350
rect 276874 514226 277494 514294
rect 276874 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 277494 514226
rect 276874 514102 277494 514170
rect 276874 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 277494 514102
rect 276874 513978 277494 514046
rect 276874 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 277494 513978
rect 276874 496350 277494 513922
rect 276874 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 277494 496350
rect 276874 496226 277494 496294
rect 276874 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 277494 496226
rect 276874 496102 277494 496170
rect 276874 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 277494 496102
rect 276874 495978 277494 496046
rect 276874 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 277494 495978
rect 276874 478350 277494 495922
rect 276874 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 277494 478350
rect 276874 478226 277494 478294
rect 276874 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 277494 478226
rect 276874 478102 277494 478170
rect 276874 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 277494 478102
rect 276874 477978 277494 478046
rect 276874 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 277494 477978
rect 276874 460350 277494 477922
rect 276874 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 277494 460350
rect 276874 460226 277494 460294
rect 276874 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 277494 460226
rect 276874 460102 277494 460170
rect 276874 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 277494 460102
rect 276874 459978 277494 460046
rect 276874 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 277494 459978
rect 276874 442350 277494 459922
rect 276874 442294 276970 442350
rect 277026 442294 277094 442350
rect 277150 442294 277218 442350
rect 277274 442294 277342 442350
rect 277398 442294 277494 442350
rect 276874 442226 277494 442294
rect 276874 442170 276970 442226
rect 277026 442170 277094 442226
rect 277150 442170 277218 442226
rect 277274 442170 277342 442226
rect 277398 442170 277494 442226
rect 276874 442102 277494 442170
rect 276874 442046 276970 442102
rect 277026 442046 277094 442102
rect 277150 442046 277218 442102
rect 277274 442046 277342 442102
rect 277398 442046 277494 442102
rect 276874 441978 277494 442046
rect 276874 441922 276970 441978
rect 277026 441922 277094 441978
rect 277150 441922 277218 441978
rect 277274 441922 277342 441978
rect 277398 441922 277494 441978
rect 276874 436006 277494 441922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 526350 291774 543922
rect 291154 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 291774 526350
rect 291154 526226 291774 526294
rect 291154 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 291774 526226
rect 291154 526102 291774 526170
rect 291154 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 291774 526102
rect 291154 525978 291774 526046
rect 291154 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 291774 525978
rect 291154 508350 291774 525922
rect 291154 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 291774 508350
rect 291154 508226 291774 508294
rect 291154 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 291774 508226
rect 291154 508102 291774 508170
rect 291154 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 291774 508102
rect 291154 507978 291774 508046
rect 291154 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 291774 507978
rect 291154 490350 291774 507922
rect 291154 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 291774 490350
rect 291154 490226 291774 490294
rect 291154 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 291774 490226
rect 291154 490102 291774 490170
rect 291154 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 291774 490102
rect 291154 489978 291774 490046
rect 291154 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 291774 489978
rect 291154 472350 291774 489922
rect 291154 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 291774 472350
rect 291154 472226 291774 472294
rect 291154 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 291774 472226
rect 291154 472102 291774 472170
rect 291154 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 291774 472102
rect 291154 471978 291774 472046
rect 291154 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 291774 471978
rect 291154 454350 291774 471922
rect 291154 454294 291250 454350
rect 291306 454294 291374 454350
rect 291430 454294 291498 454350
rect 291554 454294 291622 454350
rect 291678 454294 291774 454350
rect 291154 454226 291774 454294
rect 291154 454170 291250 454226
rect 291306 454170 291374 454226
rect 291430 454170 291498 454226
rect 291554 454170 291622 454226
rect 291678 454170 291774 454226
rect 291154 454102 291774 454170
rect 291154 454046 291250 454102
rect 291306 454046 291374 454102
rect 291430 454046 291498 454102
rect 291554 454046 291622 454102
rect 291678 454046 291774 454102
rect 291154 453978 291774 454046
rect 291154 453922 291250 453978
rect 291306 453922 291374 453978
rect 291430 453922 291498 453978
rect 291554 453922 291622 453978
rect 291678 453922 291774 453978
rect 279488 436317 279808 436380
rect 279488 436261 279558 436317
rect 279614 436261 279682 436317
rect 279738 436261 279808 436317
rect 279488 436193 279808 436261
rect 279488 436137 279558 436193
rect 279614 436137 279682 436193
rect 279738 436137 279808 436193
rect 279488 436069 279808 436137
rect 279488 436013 279558 436069
rect 279614 436013 279682 436069
rect 279738 436013 279808 436069
rect 248768 435889 248838 435945
rect 248894 435889 248962 435945
rect 249018 435889 249088 435945
rect 248768 435826 249088 435889
rect 279488 435945 279808 436013
rect 291154 436378 291774 453922
rect 294874 598172 295494 598268
rect 294874 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 295494 598172
rect 294874 598048 295494 598116
rect 294874 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 295494 598048
rect 294874 597924 295494 597992
rect 294874 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 295494 597924
rect 294874 597800 295494 597868
rect 294874 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 295494 597800
rect 294874 586350 295494 597744
rect 294874 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 295494 586350
rect 294874 586226 295494 586294
rect 294874 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 295494 586226
rect 294874 586102 295494 586170
rect 294874 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 295494 586102
rect 294874 585978 295494 586046
rect 294874 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 295494 585978
rect 294874 568350 295494 585922
rect 294874 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 295494 568350
rect 294874 568226 295494 568294
rect 294874 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 295494 568226
rect 294874 568102 295494 568170
rect 294874 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 295494 568102
rect 294874 567978 295494 568046
rect 294874 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 295494 567978
rect 294874 550350 295494 567922
rect 294874 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 295494 550350
rect 294874 550226 295494 550294
rect 294874 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 295494 550226
rect 294874 550102 295494 550170
rect 294874 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 295494 550102
rect 294874 549978 295494 550046
rect 294874 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 295494 549978
rect 294874 532350 295494 549922
rect 294874 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 295494 532350
rect 294874 532226 295494 532294
rect 294874 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 295494 532226
rect 294874 532102 295494 532170
rect 294874 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 295494 532102
rect 294874 531978 295494 532046
rect 294874 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 295494 531978
rect 294874 514350 295494 531922
rect 294874 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 295494 514350
rect 294874 514226 295494 514294
rect 294874 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 295494 514226
rect 294874 514102 295494 514170
rect 294874 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 295494 514102
rect 294874 513978 295494 514046
rect 294874 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 295494 513978
rect 294874 496350 295494 513922
rect 294874 496294 294970 496350
rect 295026 496294 295094 496350
rect 295150 496294 295218 496350
rect 295274 496294 295342 496350
rect 295398 496294 295494 496350
rect 294874 496226 295494 496294
rect 294874 496170 294970 496226
rect 295026 496170 295094 496226
rect 295150 496170 295218 496226
rect 295274 496170 295342 496226
rect 295398 496170 295494 496226
rect 294874 496102 295494 496170
rect 294874 496046 294970 496102
rect 295026 496046 295094 496102
rect 295150 496046 295218 496102
rect 295274 496046 295342 496102
rect 295398 496046 295494 496102
rect 294874 495978 295494 496046
rect 294874 495922 294970 495978
rect 295026 495922 295094 495978
rect 295150 495922 295218 495978
rect 295274 495922 295342 495978
rect 295398 495922 295494 495978
rect 294874 478350 295494 495922
rect 294874 478294 294970 478350
rect 295026 478294 295094 478350
rect 295150 478294 295218 478350
rect 295274 478294 295342 478350
rect 295398 478294 295494 478350
rect 294874 478226 295494 478294
rect 294874 478170 294970 478226
rect 295026 478170 295094 478226
rect 295150 478170 295218 478226
rect 295274 478170 295342 478226
rect 295398 478170 295494 478226
rect 294874 478102 295494 478170
rect 294874 478046 294970 478102
rect 295026 478046 295094 478102
rect 295150 478046 295218 478102
rect 295274 478046 295342 478102
rect 295398 478046 295494 478102
rect 294874 477978 295494 478046
rect 294874 477922 294970 477978
rect 295026 477922 295094 477978
rect 295150 477922 295218 477978
rect 295274 477922 295342 477978
rect 295398 477922 295494 477978
rect 294874 460350 295494 477922
rect 294874 460294 294970 460350
rect 295026 460294 295094 460350
rect 295150 460294 295218 460350
rect 295274 460294 295342 460350
rect 295398 460294 295494 460350
rect 294874 460226 295494 460294
rect 294874 460170 294970 460226
rect 295026 460170 295094 460226
rect 295150 460170 295218 460226
rect 295274 460170 295342 460226
rect 295398 460170 295494 460226
rect 294874 460102 295494 460170
rect 294874 460046 294970 460102
rect 295026 460046 295094 460102
rect 295150 460046 295218 460102
rect 295274 460046 295342 460102
rect 295398 460046 295494 460102
rect 294874 459978 295494 460046
rect 294874 459922 294970 459978
rect 295026 459922 295094 459978
rect 295150 459922 295218 459978
rect 295274 459922 295342 459978
rect 295398 459922 295494 459978
rect 294874 442350 295494 459922
rect 294874 442294 294970 442350
rect 295026 442294 295094 442350
rect 295150 442294 295218 442350
rect 295274 442294 295342 442350
rect 295398 442294 295494 442350
rect 294874 442226 295494 442294
rect 294874 442170 294970 442226
rect 295026 442170 295094 442226
rect 295150 442170 295218 442226
rect 295274 442170 295342 442226
rect 295398 442170 295494 442226
rect 294874 442102 295494 442170
rect 294874 442046 294970 442102
rect 295026 442046 295094 442102
rect 295150 442046 295218 442102
rect 295274 442046 295342 442102
rect 295398 442046 295494 442102
rect 294874 441978 295494 442046
rect 294874 441922 294970 441978
rect 295026 441922 295094 441978
rect 295150 441922 295218 441978
rect 295274 441922 295342 441978
rect 295398 441922 295494 441978
rect 294874 438436 295494 441922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 526350 309774 543922
rect 309154 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 309774 526350
rect 309154 526226 309774 526294
rect 309154 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 309774 526226
rect 309154 526102 309774 526170
rect 309154 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 309774 526102
rect 309154 525978 309774 526046
rect 309154 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 309774 525978
rect 309154 508350 309774 525922
rect 309154 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 309774 508350
rect 309154 508226 309774 508294
rect 309154 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 309774 508226
rect 309154 508102 309774 508170
rect 309154 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 309774 508102
rect 309154 507978 309774 508046
rect 309154 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 309774 507978
rect 309154 490350 309774 507922
rect 309154 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 309774 490350
rect 309154 490226 309774 490294
rect 309154 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 309774 490226
rect 309154 490102 309774 490170
rect 309154 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 309774 490102
rect 309154 489978 309774 490046
rect 309154 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 309774 489978
rect 309154 472350 309774 489922
rect 309154 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 309774 472350
rect 309154 472226 309774 472294
rect 309154 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 309774 472226
rect 309154 472102 309774 472170
rect 309154 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 309774 472102
rect 309154 471978 309774 472046
rect 309154 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 309774 471978
rect 309154 454350 309774 471922
rect 309154 454294 309250 454350
rect 309306 454294 309374 454350
rect 309430 454294 309498 454350
rect 309554 454294 309622 454350
rect 309678 454294 309774 454350
rect 309154 454226 309774 454294
rect 309154 454170 309250 454226
rect 309306 454170 309374 454226
rect 309430 454170 309498 454226
rect 309554 454170 309622 454226
rect 309678 454170 309774 454226
rect 309154 454102 309774 454170
rect 309154 454046 309250 454102
rect 309306 454046 309374 454102
rect 309430 454046 309498 454102
rect 309554 454046 309622 454102
rect 309678 454046 309774 454102
rect 309154 453978 309774 454046
rect 309154 453922 309250 453978
rect 309306 453922 309374 453978
rect 309430 453922 309498 453978
rect 309554 453922 309622 453978
rect 309678 453922 309774 453978
rect 291154 436322 291250 436378
rect 291306 436322 291374 436378
rect 291430 436322 291498 436378
rect 291554 436322 291622 436378
rect 291678 436322 291774 436378
rect 291154 436254 291774 436322
rect 291154 436198 291250 436254
rect 291306 436198 291374 436254
rect 291430 436198 291498 436254
rect 291554 436198 291622 436254
rect 291678 436198 291774 436254
rect 291154 436130 291774 436198
rect 291154 436074 291250 436130
rect 291306 436074 291374 436130
rect 291430 436074 291498 436130
rect 291554 436074 291622 436130
rect 291678 436074 291774 436130
rect 291154 436006 291774 436074
rect 309154 436378 309774 453922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 514350 313494 531922
rect 312874 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 313494 514350
rect 312874 514226 313494 514294
rect 312874 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 313494 514226
rect 312874 514102 313494 514170
rect 312874 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 313494 514102
rect 312874 513978 313494 514046
rect 312874 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 313494 513978
rect 312874 496350 313494 513922
rect 312874 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 313494 496350
rect 312874 496226 313494 496294
rect 312874 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 313494 496226
rect 312874 496102 313494 496170
rect 312874 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 313494 496102
rect 312874 495978 313494 496046
rect 312874 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 313494 495978
rect 312874 478350 313494 495922
rect 312874 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 313494 478350
rect 312874 478226 313494 478294
rect 312874 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 313494 478226
rect 312874 478102 313494 478170
rect 312874 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 313494 478102
rect 312874 477978 313494 478046
rect 312874 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 313494 477978
rect 312874 460350 313494 477922
rect 312874 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 313494 460350
rect 312874 460226 313494 460294
rect 312874 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 313494 460226
rect 312874 460102 313494 460170
rect 312874 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 313494 460102
rect 312874 459978 313494 460046
rect 312874 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 313494 459978
rect 312874 442350 313494 459922
rect 312874 442294 312970 442350
rect 313026 442294 313094 442350
rect 313150 442294 313218 442350
rect 313274 442294 313342 442350
rect 313398 442294 313494 442350
rect 312874 442226 313494 442294
rect 312874 442170 312970 442226
rect 313026 442170 313094 442226
rect 313150 442170 313218 442226
rect 313274 442170 313342 442226
rect 313398 442170 313494 442226
rect 312874 442102 313494 442170
rect 312874 442046 312970 442102
rect 313026 442046 313094 442102
rect 313150 442046 313218 442102
rect 313274 442046 313342 442102
rect 313398 442046 313494 442102
rect 312874 441978 313494 442046
rect 312874 441922 312970 441978
rect 313026 441922 313094 441978
rect 313150 441922 313218 441978
rect 313274 441922 313342 441978
rect 313398 441922 313494 441978
rect 309154 436322 309250 436378
rect 309306 436322 309374 436378
rect 309430 436322 309498 436378
rect 309554 436322 309622 436378
rect 309678 436322 309774 436378
rect 309154 436254 309774 436322
rect 309154 436198 309250 436254
rect 309306 436198 309374 436254
rect 309430 436198 309498 436254
rect 309554 436198 309622 436254
rect 309678 436198 309774 436254
rect 309154 436130 309774 436198
rect 309154 436074 309250 436130
rect 309306 436074 309374 436130
rect 309430 436074 309498 436130
rect 309554 436074 309622 436130
rect 309678 436074 309774 436130
rect 309154 436006 309774 436074
rect 310208 436317 310528 436380
rect 310208 436261 310278 436317
rect 310334 436261 310402 436317
rect 310458 436261 310528 436317
rect 310208 436193 310528 436261
rect 310208 436137 310278 436193
rect 310334 436137 310402 436193
rect 310458 436137 310528 436193
rect 310208 436069 310528 436137
rect 310208 436013 310278 436069
rect 310334 436013 310402 436069
rect 310458 436013 310528 436069
rect 279488 435889 279558 435945
rect 279614 435889 279682 435945
rect 279738 435889 279808 435945
rect 279488 435826 279808 435889
rect 310208 435945 310528 436013
rect 312874 436006 313494 441922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 526350 327774 543922
rect 327154 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 327774 526350
rect 327154 526226 327774 526294
rect 327154 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 327774 526226
rect 327154 526102 327774 526170
rect 327154 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 327774 526102
rect 327154 525978 327774 526046
rect 327154 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 327774 525978
rect 327154 508350 327774 525922
rect 327154 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 327774 508350
rect 327154 508226 327774 508294
rect 327154 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 327774 508226
rect 327154 508102 327774 508170
rect 327154 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 327774 508102
rect 327154 507978 327774 508046
rect 327154 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 327774 507978
rect 327154 490350 327774 507922
rect 327154 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 327774 490350
rect 327154 490226 327774 490294
rect 327154 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 327774 490226
rect 327154 490102 327774 490170
rect 327154 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 327774 490102
rect 327154 489978 327774 490046
rect 327154 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 327774 489978
rect 327154 472350 327774 489922
rect 327154 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 327774 472350
rect 327154 472226 327774 472294
rect 327154 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 327774 472226
rect 327154 472102 327774 472170
rect 327154 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 327774 472102
rect 327154 471978 327774 472046
rect 327154 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 327774 471978
rect 327154 454350 327774 471922
rect 327154 454294 327250 454350
rect 327306 454294 327374 454350
rect 327430 454294 327498 454350
rect 327554 454294 327622 454350
rect 327678 454294 327774 454350
rect 327154 454226 327774 454294
rect 327154 454170 327250 454226
rect 327306 454170 327374 454226
rect 327430 454170 327498 454226
rect 327554 454170 327622 454226
rect 327678 454170 327774 454226
rect 327154 454102 327774 454170
rect 327154 454046 327250 454102
rect 327306 454046 327374 454102
rect 327430 454046 327498 454102
rect 327554 454046 327622 454102
rect 327678 454046 327774 454102
rect 327154 453978 327774 454046
rect 327154 453922 327250 453978
rect 327306 453922 327374 453978
rect 327430 453922 327498 453978
rect 327554 453922 327622 453978
rect 327678 453922 327774 453978
rect 327154 436378 327774 453922
rect 327154 436322 327250 436378
rect 327306 436322 327374 436378
rect 327430 436322 327498 436378
rect 327554 436322 327622 436378
rect 327678 436322 327774 436378
rect 327154 436254 327774 436322
rect 327154 436198 327250 436254
rect 327306 436198 327374 436254
rect 327430 436198 327498 436254
rect 327554 436198 327622 436254
rect 327678 436198 327774 436254
rect 327154 436130 327774 436198
rect 327154 436074 327250 436130
rect 327306 436074 327374 436130
rect 327430 436074 327498 436130
rect 327554 436074 327622 436130
rect 327678 436074 327774 436130
rect 327154 436006 327774 436074
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 514350 331494 531922
rect 330874 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 331494 514350
rect 330874 514226 331494 514294
rect 330874 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 331494 514226
rect 330874 514102 331494 514170
rect 330874 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 331494 514102
rect 330874 513978 331494 514046
rect 330874 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 331494 513978
rect 330874 496350 331494 513922
rect 330874 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 331494 496350
rect 330874 496226 331494 496294
rect 330874 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 331494 496226
rect 330874 496102 331494 496170
rect 330874 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 331494 496102
rect 330874 495978 331494 496046
rect 330874 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 331494 495978
rect 330874 478350 331494 495922
rect 330874 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 331494 478350
rect 330874 478226 331494 478294
rect 330874 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 331494 478226
rect 330874 478102 331494 478170
rect 330874 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 331494 478102
rect 330874 477978 331494 478046
rect 330874 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 331494 477978
rect 330874 460350 331494 477922
rect 330874 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 331494 460350
rect 330874 460226 331494 460294
rect 330874 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 331494 460226
rect 330874 460102 331494 460170
rect 330874 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 331494 460102
rect 330874 459978 331494 460046
rect 330874 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 331494 459978
rect 330874 442350 331494 459922
rect 330874 442294 330970 442350
rect 331026 442294 331094 442350
rect 331150 442294 331218 442350
rect 331274 442294 331342 442350
rect 331398 442294 331494 442350
rect 330874 442226 331494 442294
rect 330874 442170 330970 442226
rect 331026 442170 331094 442226
rect 331150 442170 331218 442226
rect 331274 442170 331342 442226
rect 331398 442170 331494 442226
rect 330874 442102 331494 442170
rect 330874 442046 330970 442102
rect 331026 442046 331094 442102
rect 331150 442046 331218 442102
rect 331274 442046 331342 442102
rect 331398 442046 331494 442102
rect 330874 441978 331494 442046
rect 330874 441922 330970 441978
rect 331026 441922 331094 441978
rect 331150 441922 331218 441978
rect 331274 441922 331342 441978
rect 331398 441922 331494 441978
rect 330874 436006 331494 441922
rect 345154 597212 345774 598268
rect 345154 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 345774 597212
rect 345154 597088 345774 597156
rect 345154 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 345774 597088
rect 345154 596964 345774 597032
rect 345154 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 345774 596964
rect 345154 596840 345774 596908
rect 345154 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 345774 596840
rect 345154 580350 345774 596784
rect 345154 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 345774 580350
rect 345154 580226 345774 580294
rect 345154 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 345774 580226
rect 345154 580102 345774 580170
rect 345154 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 345774 580102
rect 345154 579978 345774 580046
rect 345154 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 345774 579978
rect 345154 562350 345774 579922
rect 345154 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 345774 562350
rect 345154 562226 345774 562294
rect 345154 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 345774 562226
rect 345154 562102 345774 562170
rect 345154 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 345774 562102
rect 345154 561978 345774 562046
rect 345154 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 345774 561978
rect 345154 544350 345774 561922
rect 345154 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 345774 544350
rect 345154 544226 345774 544294
rect 345154 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 345774 544226
rect 345154 544102 345774 544170
rect 345154 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 345774 544102
rect 345154 543978 345774 544046
rect 345154 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 345774 543978
rect 345154 526350 345774 543922
rect 345154 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 345774 526350
rect 345154 526226 345774 526294
rect 345154 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 345774 526226
rect 345154 526102 345774 526170
rect 345154 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 345774 526102
rect 345154 525978 345774 526046
rect 345154 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 345774 525978
rect 345154 508350 345774 525922
rect 345154 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 345774 508350
rect 345154 508226 345774 508294
rect 345154 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 345774 508226
rect 345154 508102 345774 508170
rect 345154 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 345774 508102
rect 345154 507978 345774 508046
rect 345154 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 345774 507978
rect 345154 490350 345774 507922
rect 345154 490294 345250 490350
rect 345306 490294 345374 490350
rect 345430 490294 345498 490350
rect 345554 490294 345622 490350
rect 345678 490294 345774 490350
rect 345154 490226 345774 490294
rect 345154 490170 345250 490226
rect 345306 490170 345374 490226
rect 345430 490170 345498 490226
rect 345554 490170 345622 490226
rect 345678 490170 345774 490226
rect 345154 490102 345774 490170
rect 345154 490046 345250 490102
rect 345306 490046 345374 490102
rect 345430 490046 345498 490102
rect 345554 490046 345622 490102
rect 345678 490046 345774 490102
rect 345154 489978 345774 490046
rect 345154 489922 345250 489978
rect 345306 489922 345374 489978
rect 345430 489922 345498 489978
rect 345554 489922 345622 489978
rect 345678 489922 345774 489978
rect 345154 472350 345774 489922
rect 345154 472294 345250 472350
rect 345306 472294 345374 472350
rect 345430 472294 345498 472350
rect 345554 472294 345622 472350
rect 345678 472294 345774 472350
rect 345154 472226 345774 472294
rect 345154 472170 345250 472226
rect 345306 472170 345374 472226
rect 345430 472170 345498 472226
rect 345554 472170 345622 472226
rect 345678 472170 345774 472226
rect 345154 472102 345774 472170
rect 345154 472046 345250 472102
rect 345306 472046 345374 472102
rect 345430 472046 345498 472102
rect 345554 472046 345622 472102
rect 345678 472046 345774 472102
rect 345154 471978 345774 472046
rect 345154 471922 345250 471978
rect 345306 471922 345374 471978
rect 345430 471922 345498 471978
rect 345554 471922 345622 471978
rect 345678 471922 345774 471978
rect 345154 454350 345774 471922
rect 345154 454294 345250 454350
rect 345306 454294 345374 454350
rect 345430 454294 345498 454350
rect 345554 454294 345622 454350
rect 345678 454294 345774 454350
rect 345154 454226 345774 454294
rect 345154 454170 345250 454226
rect 345306 454170 345374 454226
rect 345430 454170 345498 454226
rect 345554 454170 345622 454226
rect 345678 454170 345774 454226
rect 345154 454102 345774 454170
rect 345154 454046 345250 454102
rect 345306 454046 345374 454102
rect 345430 454046 345498 454102
rect 345554 454046 345622 454102
rect 345678 454046 345774 454102
rect 345154 453978 345774 454046
rect 345154 453922 345250 453978
rect 345306 453922 345374 453978
rect 345430 453922 345498 453978
rect 345554 453922 345622 453978
rect 345678 453922 345774 453978
rect 340928 436317 341248 436380
rect 340928 436261 340998 436317
rect 341054 436261 341122 436317
rect 341178 436261 341248 436317
rect 340928 436193 341248 436261
rect 340928 436137 340998 436193
rect 341054 436137 341122 436193
rect 341178 436137 341248 436193
rect 340928 436069 341248 436137
rect 340928 436013 340998 436069
rect 341054 436013 341122 436069
rect 341178 436013 341248 436069
rect 310208 435889 310278 435945
rect 310334 435889 310402 435945
rect 310458 435889 310528 435945
rect 310208 435826 310528 435889
rect 340928 435945 341248 436013
rect 345154 436378 345774 453922
rect 345154 436322 345250 436378
rect 345306 436322 345374 436378
rect 345430 436322 345498 436378
rect 345554 436322 345622 436378
rect 345678 436322 345774 436378
rect 345154 436254 345774 436322
rect 345154 436198 345250 436254
rect 345306 436198 345374 436254
rect 345430 436198 345498 436254
rect 345554 436198 345622 436254
rect 345678 436198 345774 436254
rect 345154 436130 345774 436198
rect 345154 436074 345250 436130
rect 345306 436074 345374 436130
rect 345430 436074 345498 436130
rect 345554 436074 345622 436130
rect 345678 436074 345774 436130
rect 345154 436006 345774 436074
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 514350 349494 531922
rect 348874 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 349494 514350
rect 348874 514226 349494 514294
rect 348874 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 349494 514226
rect 348874 514102 349494 514170
rect 348874 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 349494 514102
rect 348874 513978 349494 514046
rect 348874 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 349494 513978
rect 348874 496350 349494 513922
rect 348874 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 349494 496350
rect 348874 496226 349494 496294
rect 348874 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 349494 496226
rect 348874 496102 349494 496170
rect 348874 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 349494 496102
rect 348874 495978 349494 496046
rect 348874 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 349494 495978
rect 348874 478350 349494 495922
rect 348874 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 349494 478350
rect 348874 478226 349494 478294
rect 348874 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 349494 478226
rect 348874 478102 349494 478170
rect 348874 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 349494 478102
rect 348874 477978 349494 478046
rect 348874 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 349494 477978
rect 348874 460350 349494 477922
rect 348874 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 349494 460350
rect 348874 460226 349494 460294
rect 348874 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 349494 460226
rect 348874 460102 349494 460170
rect 348874 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 349494 460102
rect 348874 459978 349494 460046
rect 348874 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 349494 459978
rect 348874 442350 349494 459922
rect 348874 442294 348970 442350
rect 349026 442294 349094 442350
rect 349150 442294 349218 442350
rect 349274 442294 349342 442350
rect 349398 442294 349494 442350
rect 348874 442226 349494 442294
rect 348874 442170 348970 442226
rect 349026 442170 349094 442226
rect 349150 442170 349218 442226
rect 349274 442170 349342 442226
rect 349398 442170 349494 442226
rect 348874 442102 349494 442170
rect 348874 442046 348970 442102
rect 349026 442046 349094 442102
rect 349150 442046 349218 442102
rect 349274 442046 349342 442102
rect 349398 442046 349494 442102
rect 348874 441978 349494 442046
rect 348874 441922 348970 441978
rect 349026 441922 349094 441978
rect 349150 441922 349218 441978
rect 349274 441922 349342 441978
rect 349398 441922 349494 441978
rect 340928 435889 340998 435945
rect 341054 435889 341122 435945
rect 341178 435889 341248 435945
rect 340928 435826 341248 435889
rect 79808 424350 80128 424384
rect 79808 424294 79878 424350
rect 79934 424294 80002 424350
rect 80058 424294 80128 424350
rect 79808 424226 80128 424294
rect 79808 424170 79878 424226
rect 79934 424170 80002 424226
rect 80058 424170 80128 424226
rect 79808 424102 80128 424170
rect 79808 424046 79878 424102
rect 79934 424046 80002 424102
rect 80058 424046 80128 424102
rect 79808 423978 80128 424046
rect 79808 423922 79878 423978
rect 79934 423922 80002 423978
rect 80058 423922 80128 423978
rect 79808 423888 80128 423922
rect 110528 424350 110848 424384
rect 110528 424294 110598 424350
rect 110654 424294 110722 424350
rect 110778 424294 110848 424350
rect 110528 424226 110848 424294
rect 110528 424170 110598 424226
rect 110654 424170 110722 424226
rect 110778 424170 110848 424226
rect 110528 424102 110848 424170
rect 110528 424046 110598 424102
rect 110654 424046 110722 424102
rect 110778 424046 110848 424102
rect 110528 423978 110848 424046
rect 110528 423922 110598 423978
rect 110654 423922 110722 423978
rect 110778 423922 110848 423978
rect 110528 423888 110848 423922
rect 141248 424350 141568 424384
rect 141248 424294 141318 424350
rect 141374 424294 141442 424350
rect 141498 424294 141568 424350
rect 141248 424226 141568 424294
rect 141248 424170 141318 424226
rect 141374 424170 141442 424226
rect 141498 424170 141568 424226
rect 141248 424102 141568 424170
rect 141248 424046 141318 424102
rect 141374 424046 141442 424102
rect 141498 424046 141568 424102
rect 141248 423978 141568 424046
rect 141248 423922 141318 423978
rect 141374 423922 141442 423978
rect 141498 423922 141568 423978
rect 141248 423888 141568 423922
rect 171968 424350 172288 424384
rect 171968 424294 172038 424350
rect 172094 424294 172162 424350
rect 172218 424294 172288 424350
rect 171968 424226 172288 424294
rect 171968 424170 172038 424226
rect 172094 424170 172162 424226
rect 172218 424170 172288 424226
rect 171968 424102 172288 424170
rect 171968 424046 172038 424102
rect 172094 424046 172162 424102
rect 172218 424046 172288 424102
rect 171968 423978 172288 424046
rect 171968 423922 172038 423978
rect 172094 423922 172162 423978
rect 172218 423922 172288 423978
rect 171968 423888 172288 423922
rect 202688 424350 203008 424384
rect 202688 424294 202758 424350
rect 202814 424294 202882 424350
rect 202938 424294 203008 424350
rect 202688 424226 203008 424294
rect 202688 424170 202758 424226
rect 202814 424170 202882 424226
rect 202938 424170 203008 424226
rect 202688 424102 203008 424170
rect 202688 424046 202758 424102
rect 202814 424046 202882 424102
rect 202938 424046 203008 424102
rect 202688 423978 203008 424046
rect 202688 423922 202758 423978
rect 202814 423922 202882 423978
rect 202938 423922 203008 423978
rect 202688 423888 203008 423922
rect 233408 424350 233728 424384
rect 233408 424294 233478 424350
rect 233534 424294 233602 424350
rect 233658 424294 233728 424350
rect 233408 424226 233728 424294
rect 233408 424170 233478 424226
rect 233534 424170 233602 424226
rect 233658 424170 233728 424226
rect 233408 424102 233728 424170
rect 233408 424046 233478 424102
rect 233534 424046 233602 424102
rect 233658 424046 233728 424102
rect 233408 423978 233728 424046
rect 233408 423922 233478 423978
rect 233534 423922 233602 423978
rect 233658 423922 233728 423978
rect 233408 423888 233728 423922
rect 264128 424350 264448 424384
rect 264128 424294 264198 424350
rect 264254 424294 264322 424350
rect 264378 424294 264448 424350
rect 264128 424226 264448 424294
rect 264128 424170 264198 424226
rect 264254 424170 264322 424226
rect 264378 424170 264448 424226
rect 264128 424102 264448 424170
rect 264128 424046 264198 424102
rect 264254 424046 264322 424102
rect 264378 424046 264448 424102
rect 264128 423978 264448 424046
rect 264128 423922 264198 423978
rect 264254 423922 264322 423978
rect 264378 423922 264448 423978
rect 264128 423888 264448 423922
rect 294848 424350 295168 424384
rect 294848 424294 294918 424350
rect 294974 424294 295042 424350
rect 295098 424294 295168 424350
rect 294848 424226 295168 424294
rect 294848 424170 294918 424226
rect 294974 424170 295042 424226
rect 295098 424170 295168 424226
rect 294848 424102 295168 424170
rect 294848 424046 294918 424102
rect 294974 424046 295042 424102
rect 295098 424046 295168 424102
rect 294848 423978 295168 424046
rect 294848 423922 294918 423978
rect 294974 423922 295042 423978
rect 295098 423922 295168 423978
rect 294848 423888 295168 423922
rect 325568 424350 325888 424384
rect 325568 424294 325638 424350
rect 325694 424294 325762 424350
rect 325818 424294 325888 424350
rect 325568 424226 325888 424294
rect 325568 424170 325638 424226
rect 325694 424170 325762 424226
rect 325818 424170 325888 424226
rect 325568 424102 325888 424170
rect 325568 424046 325638 424102
rect 325694 424046 325762 424102
rect 325818 424046 325888 424102
rect 325568 423978 325888 424046
rect 325568 423922 325638 423978
rect 325694 423922 325762 423978
rect 325818 423922 325888 423978
rect 325568 423888 325888 423922
rect 348874 424350 349494 441922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 526350 363774 543922
rect 363154 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 363774 526350
rect 363154 526226 363774 526294
rect 363154 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 363774 526226
rect 363154 526102 363774 526170
rect 363154 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 363774 526102
rect 363154 525978 363774 526046
rect 363154 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 363774 525978
rect 363154 508350 363774 525922
rect 363154 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 363774 508350
rect 363154 508226 363774 508294
rect 363154 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 363774 508226
rect 363154 508102 363774 508170
rect 363154 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 363774 508102
rect 363154 507978 363774 508046
rect 363154 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 363774 507978
rect 363154 490350 363774 507922
rect 363154 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 363774 490350
rect 363154 490226 363774 490294
rect 363154 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 363774 490226
rect 363154 490102 363774 490170
rect 363154 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 363774 490102
rect 363154 489978 363774 490046
rect 363154 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 363774 489978
rect 363154 472350 363774 489922
rect 363154 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 363774 472350
rect 363154 472226 363774 472294
rect 363154 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 363774 472226
rect 363154 472102 363774 472170
rect 363154 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 363774 472102
rect 363154 471978 363774 472046
rect 363154 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 363774 471978
rect 363154 454350 363774 471922
rect 363154 454294 363250 454350
rect 363306 454294 363374 454350
rect 363430 454294 363498 454350
rect 363554 454294 363622 454350
rect 363678 454294 363774 454350
rect 363154 454226 363774 454294
rect 363154 454170 363250 454226
rect 363306 454170 363374 454226
rect 363430 454170 363498 454226
rect 363554 454170 363622 454226
rect 363678 454170 363774 454226
rect 363154 454102 363774 454170
rect 363154 454046 363250 454102
rect 363306 454046 363374 454102
rect 363430 454046 363498 454102
rect 363554 454046 363622 454102
rect 363678 454046 363774 454102
rect 363154 453978 363774 454046
rect 363154 453922 363250 453978
rect 363306 453922 363374 453978
rect 363430 453922 363498 453978
rect 363554 453922 363622 453978
rect 363678 453922 363774 453978
rect 363154 436350 363774 453922
rect 363154 436294 363250 436350
rect 363306 436294 363374 436350
rect 363430 436294 363498 436350
rect 363554 436294 363622 436350
rect 363678 436294 363774 436350
rect 363154 436226 363774 436294
rect 363154 436170 363250 436226
rect 363306 436170 363374 436226
rect 363430 436170 363498 436226
rect 363554 436170 363622 436226
rect 363678 436170 363774 436226
rect 363154 436102 363774 436170
rect 363154 436046 363250 436102
rect 363306 436046 363374 436102
rect 363430 436046 363498 436102
rect 363554 436046 363622 436102
rect 363678 436046 363774 436102
rect 363154 435978 363774 436046
rect 363154 435922 363250 435978
rect 363306 435922 363374 435978
rect 363430 435922 363498 435978
rect 363554 435922 363622 435978
rect 363678 435922 363774 435978
rect 348874 424294 348970 424350
rect 349026 424294 349094 424350
rect 349150 424294 349218 424350
rect 349274 424294 349342 424350
rect 349398 424294 349494 424350
rect 348874 424226 349494 424294
rect 348874 424170 348970 424226
rect 349026 424170 349094 424226
rect 349150 424170 349218 424226
rect 349274 424170 349342 424226
rect 349398 424170 349494 424226
rect 348874 424102 349494 424170
rect 348874 424046 348970 424102
rect 349026 424046 349094 424102
rect 349150 424046 349218 424102
rect 349274 424046 349342 424102
rect 349398 424046 349494 424102
rect 348874 423978 349494 424046
rect 348874 423922 348970 423978
rect 349026 423922 349094 423978
rect 349150 423922 349218 423978
rect 349274 423922 349342 423978
rect 349398 423922 349494 423978
rect 57154 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 57774 418350
rect 57154 418226 57774 418294
rect 57154 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 57774 418226
rect 57154 418102 57774 418170
rect 57154 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 57774 418102
rect 57154 417978 57774 418046
rect 57154 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 57774 417978
rect 57154 400350 57774 417922
rect 64448 418350 64768 418384
rect 64448 418294 64518 418350
rect 64574 418294 64642 418350
rect 64698 418294 64768 418350
rect 64448 418226 64768 418294
rect 64448 418170 64518 418226
rect 64574 418170 64642 418226
rect 64698 418170 64768 418226
rect 64448 418102 64768 418170
rect 64448 418046 64518 418102
rect 64574 418046 64642 418102
rect 64698 418046 64768 418102
rect 64448 417978 64768 418046
rect 64448 417922 64518 417978
rect 64574 417922 64642 417978
rect 64698 417922 64768 417978
rect 64448 417888 64768 417922
rect 95168 418350 95488 418384
rect 95168 418294 95238 418350
rect 95294 418294 95362 418350
rect 95418 418294 95488 418350
rect 95168 418226 95488 418294
rect 95168 418170 95238 418226
rect 95294 418170 95362 418226
rect 95418 418170 95488 418226
rect 95168 418102 95488 418170
rect 95168 418046 95238 418102
rect 95294 418046 95362 418102
rect 95418 418046 95488 418102
rect 95168 417978 95488 418046
rect 95168 417922 95238 417978
rect 95294 417922 95362 417978
rect 95418 417922 95488 417978
rect 95168 417888 95488 417922
rect 125888 418350 126208 418384
rect 125888 418294 125958 418350
rect 126014 418294 126082 418350
rect 126138 418294 126208 418350
rect 125888 418226 126208 418294
rect 125888 418170 125958 418226
rect 126014 418170 126082 418226
rect 126138 418170 126208 418226
rect 125888 418102 126208 418170
rect 125888 418046 125958 418102
rect 126014 418046 126082 418102
rect 126138 418046 126208 418102
rect 125888 417978 126208 418046
rect 125888 417922 125958 417978
rect 126014 417922 126082 417978
rect 126138 417922 126208 417978
rect 125888 417888 126208 417922
rect 156608 418350 156928 418384
rect 156608 418294 156678 418350
rect 156734 418294 156802 418350
rect 156858 418294 156928 418350
rect 156608 418226 156928 418294
rect 156608 418170 156678 418226
rect 156734 418170 156802 418226
rect 156858 418170 156928 418226
rect 156608 418102 156928 418170
rect 156608 418046 156678 418102
rect 156734 418046 156802 418102
rect 156858 418046 156928 418102
rect 156608 417978 156928 418046
rect 156608 417922 156678 417978
rect 156734 417922 156802 417978
rect 156858 417922 156928 417978
rect 156608 417888 156928 417922
rect 187328 418350 187648 418384
rect 187328 418294 187398 418350
rect 187454 418294 187522 418350
rect 187578 418294 187648 418350
rect 187328 418226 187648 418294
rect 187328 418170 187398 418226
rect 187454 418170 187522 418226
rect 187578 418170 187648 418226
rect 187328 418102 187648 418170
rect 187328 418046 187398 418102
rect 187454 418046 187522 418102
rect 187578 418046 187648 418102
rect 187328 417978 187648 418046
rect 187328 417922 187398 417978
rect 187454 417922 187522 417978
rect 187578 417922 187648 417978
rect 187328 417888 187648 417922
rect 218048 418350 218368 418384
rect 218048 418294 218118 418350
rect 218174 418294 218242 418350
rect 218298 418294 218368 418350
rect 218048 418226 218368 418294
rect 218048 418170 218118 418226
rect 218174 418170 218242 418226
rect 218298 418170 218368 418226
rect 218048 418102 218368 418170
rect 218048 418046 218118 418102
rect 218174 418046 218242 418102
rect 218298 418046 218368 418102
rect 218048 417978 218368 418046
rect 218048 417922 218118 417978
rect 218174 417922 218242 417978
rect 218298 417922 218368 417978
rect 218048 417888 218368 417922
rect 248768 418350 249088 418384
rect 248768 418294 248838 418350
rect 248894 418294 248962 418350
rect 249018 418294 249088 418350
rect 248768 418226 249088 418294
rect 248768 418170 248838 418226
rect 248894 418170 248962 418226
rect 249018 418170 249088 418226
rect 248768 418102 249088 418170
rect 248768 418046 248838 418102
rect 248894 418046 248962 418102
rect 249018 418046 249088 418102
rect 248768 417978 249088 418046
rect 248768 417922 248838 417978
rect 248894 417922 248962 417978
rect 249018 417922 249088 417978
rect 248768 417888 249088 417922
rect 279488 418350 279808 418384
rect 279488 418294 279558 418350
rect 279614 418294 279682 418350
rect 279738 418294 279808 418350
rect 279488 418226 279808 418294
rect 279488 418170 279558 418226
rect 279614 418170 279682 418226
rect 279738 418170 279808 418226
rect 279488 418102 279808 418170
rect 279488 418046 279558 418102
rect 279614 418046 279682 418102
rect 279738 418046 279808 418102
rect 279488 417978 279808 418046
rect 279488 417922 279558 417978
rect 279614 417922 279682 417978
rect 279738 417922 279808 417978
rect 279488 417888 279808 417922
rect 310208 418350 310528 418384
rect 310208 418294 310278 418350
rect 310334 418294 310402 418350
rect 310458 418294 310528 418350
rect 310208 418226 310528 418294
rect 310208 418170 310278 418226
rect 310334 418170 310402 418226
rect 310458 418170 310528 418226
rect 310208 418102 310528 418170
rect 310208 418046 310278 418102
rect 310334 418046 310402 418102
rect 310458 418046 310528 418102
rect 310208 417978 310528 418046
rect 310208 417922 310278 417978
rect 310334 417922 310402 417978
rect 310458 417922 310528 417978
rect 310208 417888 310528 417922
rect 340928 418350 341248 418384
rect 340928 418294 340998 418350
rect 341054 418294 341122 418350
rect 341178 418294 341248 418350
rect 340928 418226 341248 418294
rect 340928 418170 340998 418226
rect 341054 418170 341122 418226
rect 341178 418170 341248 418226
rect 340928 418102 341248 418170
rect 340928 418046 340998 418102
rect 341054 418046 341122 418102
rect 341178 418046 341248 418102
rect 340928 417978 341248 418046
rect 340928 417922 340998 417978
rect 341054 417922 341122 417978
rect 341178 417922 341248 417978
rect 340928 417888 341248 417922
rect 79808 406350 80128 406384
rect 79808 406294 79878 406350
rect 79934 406294 80002 406350
rect 80058 406294 80128 406350
rect 79808 406226 80128 406294
rect 79808 406170 79878 406226
rect 79934 406170 80002 406226
rect 80058 406170 80128 406226
rect 79808 406102 80128 406170
rect 79808 406046 79878 406102
rect 79934 406046 80002 406102
rect 80058 406046 80128 406102
rect 79808 405978 80128 406046
rect 79808 405922 79878 405978
rect 79934 405922 80002 405978
rect 80058 405922 80128 405978
rect 79808 405888 80128 405922
rect 110528 406350 110848 406384
rect 110528 406294 110598 406350
rect 110654 406294 110722 406350
rect 110778 406294 110848 406350
rect 110528 406226 110848 406294
rect 110528 406170 110598 406226
rect 110654 406170 110722 406226
rect 110778 406170 110848 406226
rect 110528 406102 110848 406170
rect 110528 406046 110598 406102
rect 110654 406046 110722 406102
rect 110778 406046 110848 406102
rect 110528 405978 110848 406046
rect 110528 405922 110598 405978
rect 110654 405922 110722 405978
rect 110778 405922 110848 405978
rect 110528 405888 110848 405922
rect 141248 406350 141568 406384
rect 141248 406294 141318 406350
rect 141374 406294 141442 406350
rect 141498 406294 141568 406350
rect 141248 406226 141568 406294
rect 141248 406170 141318 406226
rect 141374 406170 141442 406226
rect 141498 406170 141568 406226
rect 141248 406102 141568 406170
rect 141248 406046 141318 406102
rect 141374 406046 141442 406102
rect 141498 406046 141568 406102
rect 141248 405978 141568 406046
rect 141248 405922 141318 405978
rect 141374 405922 141442 405978
rect 141498 405922 141568 405978
rect 141248 405888 141568 405922
rect 171968 406350 172288 406384
rect 171968 406294 172038 406350
rect 172094 406294 172162 406350
rect 172218 406294 172288 406350
rect 171968 406226 172288 406294
rect 171968 406170 172038 406226
rect 172094 406170 172162 406226
rect 172218 406170 172288 406226
rect 171968 406102 172288 406170
rect 171968 406046 172038 406102
rect 172094 406046 172162 406102
rect 172218 406046 172288 406102
rect 171968 405978 172288 406046
rect 171968 405922 172038 405978
rect 172094 405922 172162 405978
rect 172218 405922 172288 405978
rect 171968 405888 172288 405922
rect 202688 406350 203008 406384
rect 202688 406294 202758 406350
rect 202814 406294 202882 406350
rect 202938 406294 203008 406350
rect 202688 406226 203008 406294
rect 202688 406170 202758 406226
rect 202814 406170 202882 406226
rect 202938 406170 203008 406226
rect 202688 406102 203008 406170
rect 202688 406046 202758 406102
rect 202814 406046 202882 406102
rect 202938 406046 203008 406102
rect 202688 405978 203008 406046
rect 202688 405922 202758 405978
rect 202814 405922 202882 405978
rect 202938 405922 203008 405978
rect 202688 405888 203008 405922
rect 233408 406350 233728 406384
rect 233408 406294 233478 406350
rect 233534 406294 233602 406350
rect 233658 406294 233728 406350
rect 233408 406226 233728 406294
rect 233408 406170 233478 406226
rect 233534 406170 233602 406226
rect 233658 406170 233728 406226
rect 233408 406102 233728 406170
rect 233408 406046 233478 406102
rect 233534 406046 233602 406102
rect 233658 406046 233728 406102
rect 233408 405978 233728 406046
rect 233408 405922 233478 405978
rect 233534 405922 233602 405978
rect 233658 405922 233728 405978
rect 233408 405888 233728 405922
rect 264128 406350 264448 406384
rect 264128 406294 264198 406350
rect 264254 406294 264322 406350
rect 264378 406294 264448 406350
rect 264128 406226 264448 406294
rect 264128 406170 264198 406226
rect 264254 406170 264322 406226
rect 264378 406170 264448 406226
rect 264128 406102 264448 406170
rect 264128 406046 264198 406102
rect 264254 406046 264322 406102
rect 264378 406046 264448 406102
rect 264128 405978 264448 406046
rect 264128 405922 264198 405978
rect 264254 405922 264322 405978
rect 264378 405922 264448 405978
rect 264128 405888 264448 405922
rect 294848 406350 295168 406384
rect 294848 406294 294918 406350
rect 294974 406294 295042 406350
rect 295098 406294 295168 406350
rect 294848 406226 295168 406294
rect 294848 406170 294918 406226
rect 294974 406170 295042 406226
rect 295098 406170 295168 406226
rect 294848 406102 295168 406170
rect 294848 406046 294918 406102
rect 294974 406046 295042 406102
rect 295098 406046 295168 406102
rect 294848 405978 295168 406046
rect 294848 405922 294918 405978
rect 294974 405922 295042 405978
rect 295098 405922 295168 405978
rect 294848 405888 295168 405922
rect 325568 406350 325888 406384
rect 325568 406294 325638 406350
rect 325694 406294 325762 406350
rect 325818 406294 325888 406350
rect 325568 406226 325888 406294
rect 325568 406170 325638 406226
rect 325694 406170 325762 406226
rect 325818 406170 325888 406226
rect 325568 406102 325888 406170
rect 325568 406046 325638 406102
rect 325694 406046 325762 406102
rect 325818 406046 325888 406102
rect 325568 405978 325888 406046
rect 325568 405922 325638 405978
rect 325694 405922 325762 405978
rect 325818 405922 325888 405978
rect 325568 405888 325888 405922
rect 348874 406350 349494 423922
rect 356288 424350 356608 424384
rect 356288 424294 356358 424350
rect 356414 424294 356482 424350
rect 356538 424294 356608 424350
rect 356288 424226 356608 424294
rect 356288 424170 356358 424226
rect 356414 424170 356482 424226
rect 356538 424170 356608 424226
rect 356288 424102 356608 424170
rect 356288 424046 356358 424102
rect 356414 424046 356482 424102
rect 356538 424046 356608 424102
rect 356288 423978 356608 424046
rect 356288 423922 356358 423978
rect 356414 423922 356482 423978
rect 356538 423922 356608 423978
rect 356288 423888 356608 423922
rect 363154 418350 363774 435922
rect 363154 418294 363250 418350
rect 363306 418294 363374 418350
rect 363430 418294 363498 418350
rect 363554 418294 363622 418350
rect 363678 418294 363774 418350
rect 363154 418226 363774 418294
rect 363154 418170 363250 418226
rect 363306 418170 363374 418226
rect 363430 418170 363498 418226
rect 363554 418170 363622 418226
rect 363678 418170 363774 418226
rect 363154 418102 363774 418170
rect 363154 418046 363250 418102
rect 363306 418046 363374 418102
rect 363430 418046 363498 418102
rect 363554 418046 363622 418102
rect 363678 418046 363774 418102
rect 363154 417978 363774 418046
rect 363154 417922 363250 417978
rect 363306 417922 363374 417978
rect 363430 417922 363498 417978
rect 363554 417922 363622 417978
rect 363678 417922 363774 417978
rect 348874 406294 348970 406350
rect 349026 406294 349094 406350
rect 349150 406294 349218 406350
rect 349274 406294 349342 406350
rect 349398 406294 349494 406350
rect 348874 406226 349494 406294
rect 348874 406170 348970 406226
rect 349026 406170 349094 406226
rect 349150 406170 349218 406226
rect 349274 406170 349342 406226
rect 349398 406170 349494 406226
rect 348874 406102 349494 406170
rect 348874 406046 348970 406102
rect 349026 406046 349094 406102
rect 349150 406046 349218 406102
rect 349274 406046 349342 406102
rect 349398 406046 349494 406102
rect 348874 405978 349494 406046
rect 348874 405922 348970 405978
rect 349026 405922 349094 405978
rect 349150 405922 349218 405978
rect 349274 405922 349342 405978
rect 349398 405922 349494 405978
rect 57154 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 57774 400350
rect 57154 400226 57774 400294
rect 57154 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 57774 400226
rect 57154 400102 57774 400170
rect 57154 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 57774 400102
rect 57154 399978 57774 400046
rect 57154 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 57774 399978
rect 57154 382350 57774 399922
rect 64448 400350 64768 400384
rect 64448 400294 64518 400350
rect 64574 400294 64642 400350
rect 64698 400294 64768 400350
rect 64448 400226 64768 400294
rect 64448 400170 64518 400226
rect 64574 400170 64642 400226
rect 64698 400170 64768 400226
rect 64448 400102 64768 400170
rect 64448 400046 64518 400102
rect 64574 400046 64642 400102
rect 64698 400046 64768 400102
rect 64448 399978 64768 400046
rect 64448 399922 64518 399978
rect 64574 399922 64642 399978
rect 64698 399922 64768 399978
rect 64448 399888 64768 399922
rect 95168 400350 95488 400384
rect 95168 400294 95238 400350
rect 95294 400294 95362 400350
rect 95418 400294 95488 400350
rect 95168 400226 95488 400294
rect 95168 400170 95238 400226
rect 95294 400170 95362 400226
rect 95418 400170 95488 400226
rect 95168 400102 95488 400170
rect 95168 400046 95238 400102
rect 95294 400046 95362 400102
rect 95418 400046 95488 400102
rect 95168 399978 95488 400046
rect 95168 399922 95238 399978
rect 95294 399922 95362 399978
rect 95418 399922 95488 399978
rect 95168 399888 95488 399922
rect 125888 400350 126208 400384
rect 125888 400294 125958 400350
rect 126014 400294 126082 400350
rect 126138 400294 126208 400350
rect 125888 400226 126208 400294
rect 125888 400170 125958 400226
rect 126014 400170 126082 400226
rect 126138 400170 126208 400226
rect 125888 400102 126208 400170
rect 125888 400046 125958 400102
rect 126014 400046 126082 400102
rect 126138 400046 126208 400102
rect 125888 399978 126208 400046
rect 125888 399922 125958 399978
rect 126014 399922 126082 399978
rect 126138 399922 126208 399978
rect 125888 399888 126208 399922
rect 156608 400350 156928 400384
rect 156608 400294 156678 400350
rect 156734 400294 156802 400350
rect 156858 400294 156928 400350
rect 156608 400226 156928 400294
rect 156608 400170 156678 400226
rect 156734 400170 156802 400226
rect 156858 400170 156928 400226
rect 156608 400102 156928 400170
rect 156608 400046 156678 400102
rect 156734 400046 156802 400102
rect 156858 400046 156928 400102
rect 156608 399978 156928 400046
rect 156608 399922 156678 399978
rect 156734 399922 156802 399978
rect 156858 399922 156928 399978
rect 156608 399888 156928 399922
rect 187328 400350 187648 400384
rect 187328 400294 187398 400350
rect 187454 400294 187522 400350
rect 187578 400294 187648 400350
rect 187328 400226 187648 400294
rect 187328 400170 187398 400226
rect 187454 400170 187522 400226
rect 187578 400170 187648 400226
rect 187328 400102 187648 400170
rect 187328 400046 187398 400102
rect 187454 400046 187522 400102
rect 187578 400046 187648 400102
rect 187328 399978 187648 400046
rect 187328 399922 187398 399978
rect 187454 399922 187522 399978
rect 187578 399922 187648 399978
rect 187328 399888 187648 399922
rect 218048 400350 218368 400384
rect 218048 400294 218118 400350
rect 218174 400294 218242 400350
rect 218298 400294 218368 400350
rect 218048 400226 218368 400294
rect 218048 400170 218118 400226
rect 218174 400170 218242 400226
rect 218298 400170 218368 400226
rect 218048 400102 218368 400170
rect 218048 400046 218118 400102
rect 218174 400046 218242 400102
rect 218298 400046 218368 400102
rect 218048 399978 218368 400046
rect 218048 399922 218118 399978
rect 218174 399922 218242 399978
rect 218298 399922 218368 399978
rect 218048 399888 218368 399922
rect 248768 400350 249088 400384
rect 248768 400294 248838 400350
rect 248894 400294 248962 400350
rect 249018 400294 249088 400350
rect 248768 400226 249088 400294
rect 248768 400170 248838 400226
rect 248894 400170 248962 400226
rect 249018 400170 249088 400226
rect 248768 400102 249088 400170
rect 248768 400046 248838 400102
rect 248894 400046 248962 400102
rect 249018 400046 249088 400102
rect 248768 399978 249088 400046
rect 248768 399922 248838 399978
rect 248894 399922 248962 399978
rect 249018 399922 249088 399978
rect 248768 399888 249088 399922
rect 279488 400350 279808 400384
rect 279488 400294 279558 400350
rect 279614 400294 279682 400350
rect 279738 400294 279808 400350
rect 279488 400226 279808 400294
rect 279488 400170 279558 400226
rect 279614 400170 279682 400226
rect 279738 400170 279808 400226
rect 279488 400102 279808 400170
rect 279488 400046 279558 400102
rect 279614 400046 279682 400102
rect 279738 400046 279808 400102
rect 279488 399978 279808 400046
rect 279488 399922 279558 399978
rect 279614 399922 279682 399978
rect 279738 399922 279808 399978
rect 279488 399888 279808 399922
rect 310208 400350 310528 400384
rect 310208 400294 310278 400350
rect 310334 400294 310402 400350
rect 310458 400294 310528 400350
rect 310208 400226 310528 400294
rect 310208 400170 310278 400226
rect 310334 400170 310402 400226
rect 310458 400170 310528 400226
rect 310208 400102 310528 400170
rect 310208 400046 310278 400102
rect 310334 400046 310402 400102
rect 310458 400046 310528 400102
rect 310208 399978 310528 400046
rect 310208 399922 310278 399978
rect 310334 399922 310402 399978
rect 310458 399922 310528 399978
rect 310208 399888 310528 399922
rect 340928 400350 341248 400384
rect 340928 400294 340998 400350
rect 341054 400294 341122 400350
rect 341178 400294 341248 400350
rect 340928 400226 341248 400294
rect 340928 400170 340998 400226
rect 341054 400170 341122 400226
rect 341178 400170 341248 400226
rect 340928 400102 341248 400170
rect 340928 400046 340998 400102
rect 341054 400046 341122 400102
rect 341178 400046 341248 400102
rect 340928 399978 341248 400046
rect 340928 399922 340998 399978
rect 341054 399922 341122 399978
rect 341178 399922 341248 399978
rect 340928 399888 341248 399922
rect 79808 388350 80128 388384
rect 79808 388294 79878 388350
rect 79934 388294 80002 388350
rect 80058 388294 80128 388350
rect 79808 388226 80128 388294
rect 79808 388170 79878 388226
rect 79934 388170 80002 388226
rect 80058 388170 80128 388226
rect 79808 388102 80128 388170
rect 79808 388046 79878 388102
rect 79934 388046 80002 388102
rect 80058 388046 80128 388102
rect 79808 387978 80128 388046
rect 79808 387922 79878 387978
rect 79934 387922 80002 387978
rect 80058 387922 80128 387978
rect 79808 387888 80128 387922
rect 110528 388350 110848 388384
rect 110528 388294 110598 388350
rect 110654 388294 110722 388350
rect 110778 388294 110848 388350
rect 110528 388226 110848 388294
rect 110528 388170 110598 388226
rect 110654 388170 110722 388226
rect 110778 388170 110848 388226
rect 110528 388102 110848 388170
rect 110528 388046 110598 388102
rect 110654 388046 110722 388102
rect 110778 388046 110848 388102
rect 110528 387978 110848 388046
rect 110528 387922 110598 387978
rect 110654 387922 110722 387978
rect 110778 387922 110848 387978
rect 110528 387888 110848 387922
rect 141248 388350 141568 388384
rect 141248 388294 141318 388350
rect 141374 388294 141442 388350
rect 141498 388294 141568 388350
rect 141248 388226 141568 388294
rect 141248 388170 141318 388226
rect 141374 388170 141442 388226
rect 141498 388170 141568 388226
rect 141248 388102 141568 388170
rect 141248 388046 141318 388102
rect 141374 388046 141442 388102
rect 141498 388046 141568 388102
rect 141248 387978 141568 388046
rect 141248 387922 141318 387978
rect 141374 387922 141442 387978
rect 141498 387922 141568 387978
rect 141248 387888 141568 387922
rect 171968 388350 172288 388384
rect 171968 388294 172038 388350
rect 172094 388294 172162 388350
rect 172218 388294 172288 388350
rect 171968 388226 172288 388294
rect 171968 388170 172038 388226
rect 172094 388170 172162 388226
rect 172218 388170 172288 388226
rect 171968 388102 172288 388170
rect 171968 388046 172038 388102
rect 172094 388046 172162 388102
rect 172218 388046 172288 388102
rect 171968 387978 172288 388046
rect 171968 387922 172038 387978
rect 172094 387922 172162 387978
rect 172218 387922 172288 387978
rect 171968 387888 172288 387922
rect 202688 388350 203008 388384
rect 202688 388294 202758 388350
rect 202814 388294 202882 388350
rect 202938 388294 203008 388350
rect 202688 388226 203008 388294
rect 202688 388170 202758 388226
rect 202814 388170 202882 388226
rect 202938 388170 203008 388226
rect 202688 388102 203008 388170
rect 202688 388046 202758 388102
rect 202814 388046 202882 388102
rect 202938 388046 203008 388102
rect 202688 387978 203008 388046
rect 202688 387922 202758 387978
rect 202814 387922 202882 387978
rect 202938 387922 203008 387978
rect 202688 387888 203008 387922
rect 233408 388350 233728 388384
rect 233408 388294 233478 388350
rect 233534 388294 233602 388350
rect 233658 388294 233728 388350
rect 233408 388226 233728 388294
rect 233408 388170 233478 388226
rect 233534 388170 233602 388226
rect 233658 388170 233728 388226
rect 233408 388102 233728 388170
rect 233408 388046 233478 388102
rect 233534 388046 233602 388102
rect 233658 388046 233728 388102
rect 233408 387978 233728 388046
rect 233408 387922 233478 387978
rect 233534 387922 233602 387978
rect 233658 387922 233728 387978
rect 233408 387888 233728 387922
rect 264128 388350 264448 388384
rect 264128 388294 264198 388350
rect 264254 388294 264322 388350
rect 264378 388294 264448 388350
rect 264128 388226 264448 388294
rect 264128 388170 264198 388226
rect 264254 388170 264322 388226
rect 264378 388170 264448 388226
rect 264128 388102 264448 388170
rect 264128 388046 264198 388102
rect 264254 388046 264322 388102
rect 264378 388046 264448 388102
rect 264128 387978 264448 388046
rect 264128 387922 264198 387978
rect 264254 387922 264322 387978
rect 264378 387922 264448 387978
rect 264128 387888 264448 387922
rect 294848 388350 295168 388384
rect 294848 388294 294918 388350
rect 294974 388294 295042 388350
rect 295098 388294 295168 388350
rect 294848 388226 295168 388294
rect 294848 388170 294918 388226
rect 294974 388170 295042 388226
rect 295098 388170 295168 388226
rect 294848 388102 295168 388170
rect 294848 388046 294918 388102
rect 294974 388046 295042 388102
rect 295098 388046 295168 388102
rect 294848 387978 295168 388046
rect 294848 387922 294918 387978
rect 294974 387922 295042 387978
rect 295098 387922 295168 387978
rect 294848 387888 295168 387922
rect 325568 388350 325888 388384
rect 325568 388294 325638 388350
rect 325694 388294 325762 388350
rect 325818 388294 325888 388350
rect 325568 388226 325888 388294
rect 325568 388170 325638 388226
rect 325694 388170 325762 388226
rect 325818 388170 325888 388226
rect 325568 388102 325888 388170
rect 325568 388046 325638 388102
rect 325694 388046 325762 388102
rect 325818 388046 325888 388102
rect 325568 387978 325888 388046
rect 325568 387922 325638 387978
rect 325694 387922 325762 387978
rect 325818 387922 325888 387978
rect 325568 387888 325888 387922
rect 348874 388350 349494 405922
rect 356288 406350 356608 406384
rect 356288 406294 356358 406350
rect 356414 406294 356482 406350
rect 356538 406294 356608 406350
rect 356288 406226 356608 406294
rect 356288 406170 356358 406226
rect 356414 406170 356482 406226
rect 356538 406170 356608 406226
rect 356288 406102 356608 406170
rect 356288 406046 356358 406102
rect 356414 406046 356482 406102
rect 356538 406046 356608 406102
rect 356288 405978 356608 406046
rect 356288 405922 356358 405978
rect 356414 405922 356482 405978
rect 356538 405922 356608 405978
rect 356288 405888 356608 405922
rect 363154 400350 363774 417922
rect 363154 400294 363250 400350
rect 363306 400294 363374 400350
rect 363430 400294 363498 400350
rect 363554 400294 363622 400350
rect 363678 400294 363774 400350
rect 363154 400226 363774 400294
rect 363154 400170 363250 400226
rect 363306 400170 363374 400226
rect 363430 400170 363498 400226
rect 363554 400170 363622 400226
rect 363678 400170 363774 400226
rect 363154 400102 363774 400170
rect 363154 400046 363250 400102
rect 363306 400046 363374 400102
rect 363430 400046 363498 400102
rect 363554 400046 363622 400102
rect 363678 400046 363774 400102
rect 363154 399978 363774 400046
rect 363154 399922 363250 399978
rect 363306 399922 363374 399978
rect 363430 399922 363498 399978
rect 363554 399922 363622 399978
rect 363678 399922 363774 399978
rect 348874 388294 348970 388350
rect 349026 388294 349094 388350
rect 349150 388294 349218 388350
rect 349274 388294 349342 388350
rect 349398 388294 349494 388350
rect 348874 388226 349494 388294
rect 348874 388170 348970 388226
rect 349026 388170 349094 388226
rect 349150 388170 349218 388226
rect 349274 388170 349342 388226
rect 349398 388170 349494 388226
rect 348874 388102 349494 388170
rect 348874 388046 348970 388102
rect 349026 388046 349094 388102
rect 349150 388046 349218 388102
rect 349274 388046 349342 388102
rect 349398 388046 349494 388102
rect 348874 387978 349494 388046
rect 348874 387922 348970 387978
rect 349026 387922 349094 387978
rect 349150 387922 349218 387978
rect 349274 387922 349342 387978
rect 349398 387922 349494 387978
rect 57154 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 57774 382350
rect 57154 382226 57774 382294
rect 57154 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 57774 382226
rect 57154 382102 57774 382170
rect 57154 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 57774 382102
rect 57154 381978 57774 382046
rect 57154 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 57774 381978
rect 57154 364350 57774 381922
rect 64448 382350 64768 382384
rect 64448 382294 64518 382350
rect 64574 382294 64642 382350
rect 64698 382294 64768 382350
rect 64448 382226 64768 382294
rect 64448 382170 64518 382226
rect 64574 382170 64642 382226
rect 64698 382170 64768 382226
rect 64448 382102 64768 382170
rect 64448 382046 64518 382102
rect 64574 382046 64642 382102
rect 64698 382046 64768 382102
rect 64448 381978 64768 382046
rect 64448 381922 64518 381978
rect 64574 381922 64642 381978
rect 64698 381922 64768 381978
rect 64448 381888 64768 381922
rect 95168 382350 95488 382384
rect 95168 382294 95238 382350
rect 95294 382294 95362 382350
rect 95418 382294 95488 382350
rect 95168 382226 95488 382294
rect 95168 382170 95238 382226
rect 95294 382170 95362 382226
rect 95418 382170 95488 382226
rect 95168 382102 95488 382170
rect 95168 382046 95238 382102
rect 95294 382046 95362 382102
rect 95418 382046 95488 382102
rect 95168 381978 95488 382046
rect 95168 381922 95238 381978
rect 95294 381922 95362 381978
rect 95418 381922 95488 381978
rect 95168 381888 95488 381922
rect 125888 382350 126208 382384
rect 125888 382294 125958 382350
rect 126014 382294 126082 382350
rect 126138 382294 126208 382350
rect 125888 382226 126208 382294
rect 125888 382170 125958 382226
rect 126014 382170 126082 382226
rect 126138 382170 126208 382226
rect 125888 382102 126208 382170
rect 125888 382046 125958 382102
rect 126014 382046 126082 382102
rect 126138 382046 126208 382102
rect 125888 381978 126208 382046
rect 125888 381922 125958 381978
rect 126014 381922 126082 381978
rect 126138 381922 126208 381978
rect 125888 381888 126208 381922
rect 156608 382350 156928 382384
rect 156608 382294 156678 382350
rect 156734 382294 156802 382350
rect 156858 382294 156928 382350
rect 156608 382226 156928 382294
rect 156608 382170 156678 382226
rect 156734 382170 156802 382226
rect 156858 382170 156928 382226
rect 156608 382102 156928 382170
rect 156608 382046 156678 382102
rect 156734 382046 156802 382102
rect 156858 382046 156928 382102
rect 156608 381978 156928 382046
rect 156608 381922 156678 381978
rect 156734 381922 156802 381978
rect 156858 381922 156928 381978
rect 156608 381888 156928 381922
rect 187328 382350 187648 382384
rect 187328 382294 187398 382350
rect 187454 382294 187522 382350
rect 187578 382294 187648 382350
rect 187328 382226 187648 382294
rect 187328 382170 187398 382226
rect 187454 382170 187522 382226
rect 187578 382170 187648 382226
rect 187328 382102 187648 382170
rect 187328 382046 187398 382102
rect 187454 382046 187522 382102
rect 187578 382046 187648 382102
rect 187328 381978 187648 382046
rect 187328 381922 187398 381978
rect 187454 381922 187522 381978
rect 187578 381922 187648 381978
rect 187328 381888 187648 381922
rect 218048 382350 218368 382384
rect 218048 382294 218118 382350
rect 218174 382294 218242 382350
rect 218298 382294 218368 382350
rect 218048 382226 218368 382294
rect 218048 382170 218118 382226
rect 218174 382170 218242 382226
rect 218298 382170 218368 382226
rect 218048 382102 218368 382170
rect 218048 382046 218118 382102
rect 218174 382046 218242 382102
rect 218298 382046 218368 382102
rect 218048 381978 218368 382046
rect 218048 381922 218118 381978
rect 218174 381922 218242 381978
rect 218298 381922 218368 381978
rect 218048 381888 218368 381922
rect 248768 382350 249088 382384
rect 248768 382294 248838 382350
rect 248894 382294 248962 382350
rect 249018 382294 249088 382350
rect 248768 382226 249088 382294
rect 248768 382170 248838 382226
rect 248894 382170 248962 382226
rect 249018 382170 249088 382226
rect 248768 382102 249088 382170
rect 248768 382046 248838 382102
rect 248894 382046 248962 382102
rect 249018 382046 249088 382102
rect 248768 381978 249088 382046
rect 248768 381922 248838 381978
rect 248894 381922 248962 381978
rect 249018 381922 249088 381978
rect 248768 381888 249088 381922
rect 279488 382350 279808 382384
rect 279488 382294 279558 382350
rect 279614 382294 279682 382350
rect 279738 382294 279808 382350
rect 279488 382226 279808 382294
rect 279488 382170 279558 382226
rect 279614 382170 279682 382226
rect 279738 382170 279808 382226
rect 279488 382102 279808 382170
rect 279488 382046 279558 382102
rect 279614 382046 279682 382102
rect 279738 382046 279808 382102
rect 279488 381978 279808 382046
rect 279488 381922 279558 381978
rect 279614 381922 279682 381978
rect 279738 381922 279808 381978
rect 279488 381888 279808 381922
rect 310208 382350 310528 382384
rect 310208 382294 310278 382350
rect 310334 382294 310402 382350
rect 310458 382294 310528 382350
rect 310208 382226 310528 382294
rect 310208 382170 310278 382226
rect 310334 382170 310402 382226
rect 310458 382170 310528 382226
rect 310208 382102 310528 382170
rect 310208 382046 310278 382102
rect 310334 382046 310402 382102
rect 310458 382046 310528 382102
rect 310208 381978 310528 382046
rect 310208 381922 310278 381978
rect 310334 381922 310402 381978
rect 310458 381922 310528 381978
rect 310208 381888 310528 381922
rect 340928 382350 341248 382384
rect 340928 382294 340998 382350
rect 341054 382294 341122 382350
rect 341178 382294 341248 382350
rect 340928 382226 341248 382294
rect 340928 382170 340998 382226
rect 341054 382170 341122 382226
rect 341178 382170 341248 382226
rect 340928 382102 341248 382170
rect 340928 382046 340998 382102
rect 341054 382046 341122 382102
rect 341178 382046 341248 382102
rect 340928 381978 341248 382046
rect 340928 381922 340998 381978
rect 341054 381922 341122 381978
rect 341178 381922 341248 381978
rect 340928 381888 341248 381922
rect 79808 370350 80128 370384
rect 79808 370294 79878 370350
rect 79934 370294 80002 370350
rect 80058 370294 80128 370350
rect 79808 370226 80128 370294
rect 79808 370170 79878 370226
rect 79934 370170 80002 370226
rect 80058 370170 80128 370226
rect 79808 370102 80128 370170
rect 79808 370046 79878 370102
rect 79934 370046 80002 370102
rect 80058 370046 80128 370102
rect 79808 369978 80128 370046
rect 79808 369922 79878 369978
rect 79934 369922 80002 369978
rect 80058 369922 80128 369978
rect 79808 369888 80128 369922
rect 110528 370350 110848 370384
rect 110528 370294 110598 370350
rect 110654 370294 110722 370350
rect 110778 370294 110848 370350
rect 110528 370226 110848 370294
rect 110528 370170 110598 370226
rect 110654 370170 110722 370226
rect 110778 370170 110848 370226
rect 110528 370102 110848 370170
rect 110528 370046 110598 370102
rect 110654 370046 110722 370102
rect 110778 370046 110848 370102
rect 110528 369978 110848 370046
rect 110528 369922 110598 369978
rect 110654 369922 110722 369978
rect 110778 369922 110848 369978
rect 110528 369888 110848 369922
rect 141248 370350 141568 370384
rect 141248 370294 141318 370350
rect 141374 370294 141442 370350
rect 141498 370294 141568 370350
rect 141248 370226 141568 370294
rect 141248 370170 141318 370226
rect 141374 370170 141442 370226
rect 141498 370170 141568 370226
rect 141248 370102 141568 370170
rect 141248 370046 141318 370102
rect 141374 370046 141442 370102
rect 141498 370046 141568 370102
rect 141248 369978 141568 370046
rect 141248 369922 141318 369978
rect 141374 369922 141442 369978
rect 141498 369922 141568 369978
rect 141248 369888 141568 369922
rect 171968 370350 172288 370384
rect 171968 370294 172038 370350
rect 172094 370294 172162 370350
rect 172218 370294 172288 370350
rect 171968 370226 172288 370294
rect 171968 370170 172038 370226
rect 172094 370170 172162 370226
rect 172218 370170 172288 370226
rect 171968 370102 172288 370170
rect 171968 370046 172038 370102
rect 172094 370046 172162 370102
rect 172218 370046 172288 370102
rect 171968 369978 172288 370046
rect 171968 369922 172038 369978
rect 172094 369922 172162 369978
rect 172218 369922 172288 369978
rect 171968 369888 172288 369922
rect 202688 370350 203008 370384
rect 202688 370294 202758 370350
rect 202814 370294 202882 370350
rect 202938 370294 203008 370350
rect 202688 370226 203008 370294
rect 202688 370170 202758 370226
rect 202814 370170 202882 370226
rect 202938 370170 203008 370226
rect 202688 370102 203008 370170
rect 202688 370046 202758 370102
rect 202814 370046 202882 370102
rect 202938 370046 203008 370102
rect 202688 369978 203008 370046
rect 202688 369922 202758 369978
rect 202814 369922 202882 369978
rect 202938 369922 203008 369978
rect 202688 369888 203008 369922
rect 233408 370350 233728 370384
rect 233408 370294 233478 370350
rect 233534 370294 233602 370350
rect 233658 370294 233728 370350
rect 233408 370226 233728 370294
rect 233408 370170 233478 370226
rect 233534 370170 233602 370226
rect 233658 370170 233728 370226
rect 233408 370102 233728 370170
rect 233408 370046 233478 370102
rect 233534 370046 233602 370102
rect 233658 370046 233728 370102
rect 233408 369978 233728 370046
rect 233408 369922 233478 369978
rect 233534 369922 233602 369978
rect 233658 369922 233728 369978
rect 233408 369888 233728 369922
rect 264128 370350 264448 370384
rect 264128 370294 264198 370350
rect 264254 370294 264322 370350
rect 264378 370294 264448 370350
rect 264128 370226 264448 370294
rect 264128 370170 264198 370226
rect 264254 370170 264322 370226
rect 264378 370170 264448 370226
rect 264128 370102 264448 370170
rect 264128 370046 264198 370102
rect 264254 370046 264322 370102
rect 264378 370046 264448 370102
rect 264128 369978 264448 370046
rect 264128 369922 264198 369978
rect 264254 369922 264322 369978
rect 264378 369922 264448 369978
rect 264128 369888 264448 369922
rect 294848 370350 295168 370384
rect 294848 370294 294918 370350
rect 294974 370294 295042 370350
rect 295098 370294 295168 370350
rect 294848 370226 295168 370294
rect 294848 370170 294918 370226
rect 294974 370170 295042 370226
rect 295098 370170 295168 370226
rect 294848 370102 295168 370170
rect 294848 370046 294918 370102
rect 294974 370046 295042 370102
rect 295098 370046 295168 370102
rect 294848 369978 295168 370046
rect 294848 369922 294918 369978
rect 294974 369922 295042 369978
rect 295098 369922 295168 369978
rect 294848 369888 295168 369922
rect 325568 370350 325888 370384
rect 325568 370294 325638 370350
rect 325694 370294 325762 370350
rect 325818 370294 325888 370350
rect 325568 370226 325888 370294
rect 325568 370170 325638 370226
rect 325694 370170 325762 370226
rect 325818 370170 325888 370226
rect 325568 370102 325888 370170
rect 325568 370046 325638 370102
rect 325694 370046 325762 370102
rect 325818 370046 325888 370102
rect 325568 369978 325888 370046
rect 325568 369922 325638 369978
rect 325694 369922 325762 369978
rect 325818 369922 325888 369978
rect 325568 369888 325888 369922
rect 348874 370350 349494 387922
rect 356288 388350 356608 388384
rect 356288 388294 356358 388350
rect 356414 388294 356482 388350
rect 356538 388294 356608 388350
rect 356288 388226 356608 388294
rect 356288 388170 356358 388226
rect 356414 388170 356482 388226
rect 356538 388170 356608 388226
rect 356288 388102 356608 388170
rect 356288 388046 356358 388102
rect 356414 388046 356482 388102
rect 356538 388046 356608 388102
rect 356288 387978 356608 388046
rect 356288 387922 356358 387978
rect 356414 387922 356482 387978
rect 356538 387922 356608 387978
rect 356288 387888 356608 387922
rect 363154 382350 363774 399922
rect 363154 382294 363250 382350
rect 363306 382294 363374 382350
rect 363430 382294 363498 382350
rect 363554 382294 363622 382350
rect 363678 382294 363774 382350
rect 363154 382226 363774 382294
rect 363154 382170 363250 382226
rect 363306 382170 363374 382226
rect 363430 382170 363498 382226
rect 363554 382170 363622 382226
rect 363678 382170 363774 382226
rect 363154 382102 363774 382170
rect 363154 382046 363250 382102
rect 363306 382046 363374 382102
rect 363430 382046 363498 382102
rect 363554 382046 363622 382102
rect 363678 382046 363774 382102
rect 363154 381978 363774 382046
rect 363154 381922 363250 381978
rect 363306 381922 363374 381978
rect 363430 381922 363498 381978
rect 363554 381922 363622 381978
rect 363678 381922 363774 381978
rect 348874 370294 348970 370350
rect 349026 370294 349094 370350
rect 349150 370294 349218 370350
rect 349274 370294 349342 370350
rect 349398 370294 349494 370350
rect 348874 370226 349494 370294
rect 348874 370170 348970 370226
rect 349026 370170 349094 370226
rect 349150 370170 349218 370226
rect 349274 370170 349342 370226
rect 349398 370170 349494 370226
rect 348874 370102 349494 370170
rect 348874 370046 348970 370102
rect 349026 370046 349094 370102
rect 349150 370046 349218 370102
rect 349274 370046 349342 370102
rect 349398 370046 349494 370102
rect 348874 369978 349494 370046
rect 348874 369922 348970 369978
rect 349026 369922 349094 369978
rect 349150 369922 349218 369978
rect 349274 369922 349342 369978
rect 349398 369922 349494 369978
rect 57154 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 57774 364350
rect 57154 364226 57774 364294
rect 57154 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 57774 364226
rect 57154 364102 57774 364170
rect 57154 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 57774 364102
rect 57154 363978 57774 364046
rect 57154 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 57774 363978
rect 57154 346350 57774 363922
rect 64448 364350 64768 364384
rect 64448 364294 64518 364350
rect 64574 364294 64642 364350
rect 64698 364294 64768 364350
rect 64448 364226 64768 364294
rect 64448 364170 64518 364226
rect 64574 364170 64642 364226
rect 64698 364170 64768 364226
rect 64448 364102 64768 364170
rect 64448 364046 64518 364102
rect 64574 364046 64642 364102
rect 64698 364046 64768 364102
rect 64448 363978 64768 364046
rect 64448 363922 64518 363978
rect 64574 363922 64642 363978
rect 64698 363922 64768 363978
rect 64448 363888 64768 363922
rect 95168 364350 95488 364384
rect 95168 364294 95238 364350
rect 95294 364294 95362 364350
rect 95418 364294 95488 364350
rect 95168 364226 95488 364294
rect 95168 364170 95238 364226
rect 95294 364170 95362 364226
rect 95418 364170 95488 364226
rect 95168 364102 95488 364170
rect 95168 364046 95238 364102
rect 95294 364046 95362 364102
rect 95418 364046 95488 364102
rect 95168 363978 95488 364046
rect 95168 363922 95238 363978
rect 95294 363922 95362 363978
rect 95418 363922 95488 363978
rect 95168 363888 95488 363922
rect 125888 364350 126208 364384
rect 125888 364294 125958 364350
rect 126014 364294 126082 364350
rect 126138 364294 126208 364350
rect 125888 364226 126208 364294
rect 125888 364170 125958 364226
rect 126014 364170 126082 364226
rect 126138 364170 126208 364226
rect 125888 364102 126208 364170
rect 125888 364046 125958 364102
rect 126014 364046 126082 364102
rect 126138 364046 126208 364102
rect 125888 363978 126208 364046
rect 125888 363922 125958 363978
rect 126014 363922 126082 363978
rect 126138 363922 126208 363978
rect 125888 363888 126208 363922
rect 156608 364350 156928 364384
rect 156608 364294 156678 364350
rect 156734 364294 156802 364350
rect 156858 364294 156928 364350
rect 156608 364226 156928 364294
rect 156608 364170 156678 364226
rect 156734 364170 156802 364226
rect 156858 364170 156928 364226
rect 156608 364102 156928 364170
rect 156608 364046 156678 364102
rect 156734 364046 156802 364102
rect 156858 364046 156928 364102
rect 156608 363978 156928 364046
rect 156608 363922 156678 363978
rect 156734 363922 156802 363978
rect 156858 363922 156928 363978
rect 156608 363888 156928 363922
rect 187328 364350 187648 364384
rect 187328 364294 187398 364350
rect 187454 364294 187522 364350
rect 187578 364294 187648 364350
rect 187328 364226 187648 364294
rect 187328 364170 187398 364226
rect 187454 364170 187522 364226
rect 187578 364170 187648 364226
rect 187328 364102 187648 364170
rect 187328 364046 187398 364102
rect 187454 364046 187522 364102
rect 187578 364046 187648 364102
rect 187328 363978 187648 364046
rect 187328 363922 187398 363978
rect 187454 363922 187522 363978
rect 187578 363922 187648 363978
rect 187328 363888 187648 363922
rect 218048 364350 218368 364384
rect 218048 364294 218118 364350
rect 218174 364294 218242 364350
rect 218298 364294 218368 364350
rect 218048 364226 218368 364294
rect 218048 364170 218118 364226
rect 218174 364170 218242 364226
rect 218298 364170 218368 364226
rect 218048 364102 218368 364170
rect 218048 364046 218118 364102
rect 218174 364046 218242 364102
rect 218298 364046 218368 364102
rect 218048 363978 218368 364046
rect 218048 363922 218118 363978
rect 218174 363922 218242 363978
rect 218298 363922 218368 363978
rect 218048 363888 218368 363922
rect 248768 364350 249088 364384
rect 248768 364294 248838 364350
rect 248894 364294 248962 364350
rect 249018 364294 249088 364350
rect 248768 364226 249088 364294
rect 248768 364170 248838 364226
rect 248894 364170 248962 364226
rect 249018 364170 249088 364226
rect 248768 364102 249088 364170
rect 248768 364046 248838 364102
rect 248894 364046 248962 364102
rect 249018 364046 249088 364102
rect 248768 363978 249088 364046
rect 248768 363922 248838 363978
rect 248894 363922 248962 363978
rect 249018 363922 249088 363978
rect 248768 363888 249088 363922
rect 279488 364350 279808 364384
rect 279488 364294 279558 364350
rect 279614 364294 279682 364350
rect 279738 364294 279808 364350
rect 279488 364226 279808 364294
rect 279488 364170 279558 364226
rect 279614 364170 279682 364226
rect 279738 364170 279808 364226
rect 279488 364102 279808 364170
rect 279488 364046 279558 364102
rect 279614 364046 279682 364102
rect 279738 364046 279808 364102
rect 279488 363978 279808 364046
rect 279488 363922 279558 363978
rect 279614 363922 279682 363978
rect 279738 363922 279808 363978
rect 279488 363888 279808 363922
rect 310208 364350 310528 364384
rect 310208 364294 310278 364350
rect 310334 364294 310402 364350
rect 310458 364294 310528 364350
rect 310208 364226 310528 364294
rect 310208 364170 310278 364226
rect 310334 364170 310402 364226
rect 310458 364170 310528 364226
rect 310208 364102 310528 364170
rect 310208 364046 310278 364102
rect 310334 364046 310402 364102
rect 310458 364046 310528 364102
rect 310208 363978 310528 364046
rect 310208 363922 310278 363978
rect 310334 363922 310402 363978
rect 310458 363922 310528 363978
rect 310208 363888 310528 363922
rect 340928 364350 341248 364384
rect 340928 364294 340998 364350
rect 341054 364294 341122 364350
rect 341178 364294 341248 364350
rect 340928 364226 341248 364294
rect 340928 364170 340998 364226
rect 341054 364170 341122 364226
rect 341178 364170 341248 364226
rect 340928 364102 341248 364170
rect 340928 364046 340998 364102
rect 341054 364046 341122 364102
rect 341178 364046 341248 364102
rect 340928 363978 341248 364046
rect 340928 363922 340998 363978
rect 341054 363922 341122 363978
rect 341178 363922 341248 363978
rect 340928 363888 341248 363922
rect 79808 352350 80128 352384
rect 79808 352294 79878 352350
rect 79934 352294 80002 352350
rect 80058 352294 80128 352350
rect 79808 352226 80128 352294
rect 79808 352170 79878 352226
rect 79934 352170 80002 352226
rect 80058 352170 80128 352226
rect 79808 352102 80128 352170
rect 79808 352046 79878 352102
rect 79934 352046 80002 352102
rect 80058 352046 80128 352102
rect 79808 351978 80128 352046
rect 79808 351922 79878 351978
rect 79934 351922 80002 351978
rect 80058 351922 80128 351978
rect 79808 351888 80128 351922
rect 110528 352350 110848 352384
rect 110528 352294 110598 352350
rect 110654 352294 110722 352350
rect 110778 352294 110848 352350
rect 110528 352226 110848 352294
rect 110528 352170 110598 352226
rect 110654 352170 110722 352226
rect 110778 352170 110848 352226
rect 110528 352102 110848 352170
rect 110528 352046 110598 352102
rect 110654 352046 110722 352102
rect 110778 352046 110848 352102
rect 110528 351978 110848 352046
rect 110528 351922 110598 351978
rect 110654 351922 110722 351978
rect 110778 351922 110848 351978
rect 110528 351888 110848 351922
rect 141248 352350 141568 352384
rect 141248 352294 141318 352350
rect 141374 352294 141442 352350
rect 141498 352294 141568 352350
rect 141248 352226 141568 352294
rect 141248 352170 141318 352226
rect 141374 352170 141442 352226
rect 141498 352170 141568 352226
rect 141248 352102 141568 352170
rect 141248 352046 141318 352102
rect 141374 352046 141442 352102
rect 141498 352046 141568 352102
rect 141248 351978 141568 352046
rect 141248 351922 141318 351978
rect 141374 351922 141442 351978
rect 141498 351922 141568 351978
rect 141248 351888 141568 351922
rect 171968 352350 172288 352384
rect 171968 352294 172038 352350
rect 172094 352294 172162 352350
rect 172218 352294 172288 352350
rect 171968 352226 172288 352294
rect 171968 352170 172038 352226
rect 172094 352170 172162 352226
rect 172218 352170 172288 352226
rect 171968 352102 172288 352170
rect 171968 352046 172038 352102
rect 172094 352046 172162 352102
rect 172218 352046 172288 352102
rect 171968 351978 172288 352046
rect 171968 351922 172038 351978
rect 172094 351922 172162 351978
rect 172218 351922 172288 351978
rect 171968 351888 172288 351922
rect 202688 352350 203008 352384
rect 202688 352294 202758 352350
rect 202814 352294 202882 352350
rect 202938 352294 203008 352350
rect 202688 352226 203008 352294
rect 202688 352170 202758 352226
rect 202814 352170 202882 352226
rect 202938 352170 203008 352226
rect 202688 352102 203008 352170
rect 202688 352046 202758 352102
rect 202814 352046 202882 352102
rect 202938 352046 203008 352102
rect 202688 351978 203008 352046
rect 202688 351922 202758 351978
rect 202814 351922 202882 351978
rect 202938 351922 203008 351978
rect 202688 351888 203008 351922
rect 233408 352350 233728 352384
rect 233408 352294 233478 352350
rect 233534 352294 233602 352350
rect 233658 352294 233728 352350
rect 233408 352226 233728 352294
rect 233408 352170 233478 352226
rect 233534 352170 233602 352226
rect 233658 352170 233728 352226
rect 233408 352102 233728 352170
rect 233408 352046 233478 352102
rect 233534 352046 233602 352102
rect 233658 352046 233728 352102
rect 233408 351978 233728 352046
rect 233408 351922 233478 351978
rect 233534 351922 233602 351978
rect 233658 351922 233728 351978
rect 233408 351888 233728 351922
rect 264128 352350 264448 352384
rect 264128 352294 264198 352350
rect 264254 352294 264322 352350
rect 264378 352294 264448 352350
rect 264128 352226 264448 352294
rect 264128 352170 264198 352226
rect 264254 352170 264322 352226
rect 264378 352170 264448 352226
rect 264128 352102 264448 352170
rect 264128 352046 264198 352102
rect 264254 352046 264322 352102
rect 264378 352046 264448 352102
rect 264128 351978 264448 352046
rect 264128 351922 264198 351978
rect 264254 351922 264322 351978
rect 264378 351922 264448 351978
rect 264128 351888 264448 351922
rect 294848 352350 295168 352384
rect 294848 352294 294918 352350
rect 294974 352294 295042 352350
rect 295098 352294 295168 352350
rect 294848 352226 295168 352294
rect 294848 352170 294918 352226
rect 294974 352170 295042 352226
rect 295098 352170 295168 352226
rect 294848 352102 295168 352170
rect 294848 352046 294918 352102
rect 294974 352046 295042 352102
rect 295098 352046 295168 352102
rect 294848 351978 295168 352046
rect 294848 351922 294918 351978
rect 294974 351922 295042 351978
rect 295098 351922 295168 351978
rect 294848 351888 295168 351922
rect 325568 352350 325888 352384
rect 325568 352294 325638 352350
rect 325694 352294 325762 352350
rect 325818 352294 325888 352350
rect 325568 352226 325888 352294
rect 325568 352170 325638 352226
rect 325694 352170 325762 352226
rect 325818 352170 325888 352226
rect 325568 352102 325888 352170
rect 325568 352046 325638 352102
rect 325694 352046 325762 352102
rect 325818 352046 325888 352102
rect 325568 351978 325888 352046
rect 325568 351922 325638 351978
rect 325694 351922 325762 351978
rect 325818 351922 325888 351978
rect 325568 351888 325888 351922
rect 348874 352350 349494 369922
rect 356288 370350 356608 370384
rect 356288 370294 356358 370350
rect 356414 370294 356482 370350
rect 356538 370294 356608 370350
rect 356288 370226 356608 370294
rect 356288 370170 356358 370226
rect 356414 370170 356482 370226
rect 356538 370170 356608 370226
rect 356288 370102 356608 370170
rect 356288 370046 356358 370102
rect 356414 370046 356482 370102
rect 356538 370046 356608 370102
rect 356288 369978 356608 370046
rect 356288 369922 356358 369978
rect 356414 369922 356482 369978
rect 356538 369922 356608 369978
rect 356288 369888 356608 369922
rect 363154 364350 363774 381922
rect 363154 364294 363250 364350
rect 363306 364294 363374 364350
rect 363430 364294 363498 364350
rect 363554 364294 363622 364350
rect 363678 364294 363774 364350
rect 363154 364226 363774 364294
rect 363154 364170 363250 364226
rect 363306 364170 363374 364226
rect 363430 364170 363498 364226
rect 363554 364170 363622 364226
rect 363678 364170 363774 364226
rect 363154 364102 363774 364170
rect 363154 364046 363250 364102
rect 363306 364046 363374 364102
rect 363430 364046 363498 364102
rect 363554 364046 363622 364102
rect 363678 364046 363774 364102
rect 363154 363978 363774 364046
rect 363154 363922 363250 363978
rect 363306 363922 363374 363978
rect 363430 363922 363498 363978
rect 363554 363922 363622 363978
rect 363678 363922 363774 363978
rect 348874 352294 348970 352350
rect 349026 352294 349094 352350
rect 349150 352294 349218 352350
rect 349274 352294 349342 352350
rect 349398 352294 349494 352350
rect 348874 352226 349494 352294
rect 348874 352170 348970 352226
rect 349026 352170 349094 352226
rect 349150 352170 349218 352226
rect 349274 352170 349342 352226
rect 349398 352170 349494 352226
rect 348874 352102 349494 352170
rect 348874 352046 348970 352102
rect 349026 352046 349094 352102
rect 349150 352046 349218 352102
rect 349274 352046 349342 352102
rect 349398 352046 349494 352102
rect 348874 351978 349494 352046
rect 348874 351922 348970 351978
rect 349026 351922 349094 351978
rect 349150 351922 349218 351978
rect 349274 351922 349342 351978
rect 349398 351922 349494 351978
rect 57154 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 57774 346350
rect 57154 346226 57774 346294
rect 57154 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 57774 346226
rect 57154 346102 57774 346170
rect 57154 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 57774 346102
rect 57154 345978 57774 346046
rect 57154 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 57774 345978
rect 57154 328350 57774 345922
rect 64448 346350 64768 346384
rect 64448 346294 64518 346350
rect 64574 346294 64642 346350
rect 64698 346294 64768 346350
rect 64448 346226 64768 346294
rect 64448 346170 64518 346226
rect 64574 346170 64642 346226
rect 64698 346170 64768 346226
rect 64448 346102 64768 346170
rect 64448 346046 64518 346102
rect 64574 346046 64642 346102
rect 64698 346046 64768 346102
rect 64448 345978 64768 346046
rect 64448 345922 64518 345978
rect 64574 345922 64642 345978
rect 64698 345922 64768 345978
rect 64448 345888 64768 345922
rect 95168 346350 95488 346384
rect 95168 346294 95238 346350
rect 95294 346294 95362 346350
rect 95418 346294 95488 346350
rect 95168 346226 95488 346294
rect 95168 346170 95238 346226
rect 95294 346170 95362 346226
rect 95418 346170 95488 346226
rect 95168 346102 95488 346170
rect 95168 346046 95238 346102
rect 95294 346046 95362 346102
rect 95418 346046 95488 346102
rect 95168 345978 95488 346046
rect 95168 345922 95238 345978
rect 95294 345922 95362 345978
rect 95418 345922 95488 345978
rect 95168 345888 95488 345922
rect 125888 346350 126208 346384
rect 125888 346294 125958 346350
rect 126014 346294 126082 346350
rect 126138 346294 126208 346350
rect 125888 346226 126208 346294
rect 125888 346170 125958 346226
rect 126014 346170 126082 346226
rect 126138 346170 126208 346226
rect 125888 346102 126208 346170
rect 125888 346046 125958 346102
rect 126014 346046 126082 346102
rect 126138 346046 126208 346102
rect 125888 345978 126208 346046
rect 125888 345922 125958 345978
rect 126014 345922 126082 345978
rect 126138 345922 126208 345978
rect 125888 345888 126208 345922
rect 156608 346350 156928 346384
rect 156608 346294 156678 346350
rect 156734 346294 156802 346350
rect 156858 346294 156928 346350
rect 156608 346226 156928 346294
rect 156608 346170 156678 346226
rect 156734 346170 156802 346226
rect 156858 346170 156928 346226
rect 156608 346102 156928 346170
rect 156608 346046 156678 346102
rect 156734 346046 156802 346102
rect 156858 346046 156928 346102
rect 156608 345978 156928 346046
rect 156608 345922 156678 345978
rect 156734 345922 156802 345978
rect 156858 345922 156928 345978
rect 156608 345888 156928 345922
rect 187328 346350 187648 346384
rect 187328 346294 187398 346350
rect 187454 346294 187522 346350
rect 187578 346294 187648 346350
rect 187328 346226 187648 346294
rect 187328 346170 187398 346226
rect 187454 346170 187522 346226
rect 187578 346170 187648 346226
rect 187328 346102 187648 346170
rect 187328 346046 187398 346102
rect 187454 346046 187522 346102
rect 187578 346046 187648 346102
rect 187328 345978 187648 346046
rect 187328 345922 187398 345978
rect 187454 345922 187522 345978
rect 187578 345922 187648 345978
rect 187328 345888 187648 345922
rect 218048 346350 218368 346384
rect 218048 346294 218118 346350
rect 218174 346294 218242 346350
rect 218298 346294 218368 346350
rect 218048 346226 218368 346294
rect 218048 346170 218118 346226
rect 218174 346170 218242 346226
rect 218298 346170 218368 346226
rect 218048 346102 218368 346170
rect 218048 346046 218118 346102
rect 218174 346046 218242 346102
rect 218298 346046 218368 346102
rect 218048 345978 218368 346046
rect 218048 345922 218118 345978
rect 218174 345922 218242 345978
rect 218298 345922 218368 345978
rect 218048 345888 218368 345922
rect 248768 346350 249088 346384
rect 248768 346294 248838 346350
rect 248894 346294 248962 346350
rect 249018 346294 249088 346350
rect 248768 346226 249088 346294
rect 248768 346170 248838 346226
rect 248894 346170 248962 346226
rect 249018 346170 249088 346226
rect 248768 346102 249088 346170
rect 248768 346046 248838 346102
rect 248894 346046 248962 346102
rect 249018 346046 249088 346102
rect 248768 345978 249088 346046
rect 248768 345922 248838 345978
rect 248894 345922 248962 345978
rect 249018 345922 249088 345978
rect 248768 345888 249088 345922
rect 279488 346350 279808 346384
rect 279488 346294 279558 346350
rect 279614 346294 279682 346350
rect 279738 346294 279808 346350
rect 279488 346226 279808 346294
rect 279488 346170 279558 346226
rect 279614 346170 279682 346226
rect 279738 346170 279808 346226
rect 279488 346102 279808 346170
rect 279488 346046 279558 346102
rect 279614 346046 279682 346102
rect 279738 346046 279808 346102
rect 279488 345978 279808 346046
rect 279488 345922 279558 345978
rect 279614 345922 279682 345978
rect 279738 345922 279808 345978
rect 279488 345888 279808 345922
rect 310208 346350 310528 346384
rect 310208 346294 310278 346350
rect 310334 346294 310402 346350
rect 310458 346294 310528 346350
rect 310208 346226 310528 346294
rect 310208 346170 310278 346226
rect 310334 346170 310402 346226
rect 310458 346170 310528 346226
rect 310208 346102 310528 346170
rect 310208 346046 310278 346102
rect 310334 346046 310402 346102
rect 310458 346046 310528 346102
rect 310208 345978 310528 346046
rect 310208 345922 310278 345978
rect 310334 345922 310402 345978
rect 310458 345922 310528 345978
rect 310208 345888 310528 345922
rect 340928 346350 341248 346384
rect 340928 346294 340998 346350
rect 341054 346294 341122 346350
rect 341178 346294 341248 346350
rect 340928 346226 341248 346294
rect 340928 346170 340998 346226
rect 341054 346170 341122 346226
rect 341178 346170 341248 346226
rect 340928 346102 341248 346170
rect 340928 346046 340998 346102
rect 341054 346046 341122 346102
rect 341178 346046 341248 346102
rect 340928 345978 341248 346046
rect 340928 345922 340998 345978
rect 341054 345922 341122 345978
rect 341178 345922 341248 345978
rect 340928 345888 341248 345922
rect 79808 334350 80128 334384
rect 79808 334294 79878 334350
rect 79934 334294 80002 334350
rect 80058 334294 80128 334350
rect 79808 334226 80128 334294
rect 79808 334170 79878 334226
rect 79934 334170 80002 334226
rect 80058 334170 80128 334226
rect 79808 334102 80128 334170
rect 79808 334046 79878 334102
rect 79934 334046 80002 334102
rect 80058 334046 80128 334102
rect 79808 333978 80128 334046
rect 79808 333922 79878 333978
rect 79934 333922 80002 333978
rect 80058 333922 80128 333978
rect 79808 333888 80128 333922
rect 110528 334350 110848 334384
rect 110528 334294 110598 334350
rect 110654 334294 110722 334350
rect 110778 334294 110848 334350
rect 110528 334226 110848 334294
rect 110528 334170 110598 334226
rect 110654 334170 110722 334226
rect 110778 334170 110848 334226
rect 110528 334102 110848 334170
rect 110528 334046 110598 334102
rect 110654 334046 110722 334102
rect 110778 334046 110848 334102
rect 110528 333978 110848 334046
rect 110528 333922 110598 333978
rect 110654 333922 110722 333978
rect 110778 333922 110848 333978
rect 110528 333888 110848 333922
rect 141248 334350 141568 334384
rect 141248 334294 141318 334350
rect 141374 334294 141442 334350
rect 141498 334294 141568 334350
rect 141248 334226 141568 334294
rect 141248 334170 141318 334226
rect 141374 334170 141442 334226
rect 141498 334170 141568 334226
rect 141248 334102 141568 334170
rect 141248 334046 141318 334102
rect 141374 334046 141442 334102
rect 141498 334046 141568 334102
rect 141248 333978 141568 334046
rect 141248 333922 141318 333978
rect 141374 333922 141442 333978
rect 141498 333922 141568 333978
rect 141248 333888 141568 333922
rect 171968 334350 172288 334384
rect 171968 334294 172038 334350
rect 172094 334294 172162 334350
rect 172218 334294 172288 334350
rect 171968 334226 172288 334294
rect 171968 334170 172038 334226
rect 172094 334170 172162 334226
rect 172218 334170 172288 334226
rect 171968 334102 172288 334170
rect 171968 334046 172038 334102
rect 172094 334046 172162 334102
rect 172218 334046 172288 334102
rect 171968 333978 172288 334046
rect 171968 333922 172038 333978
rect 172094 333922 172162 333978
rect 172218 333922 172288 333978
rect 171968 333888 172288 333922
rect 202688 334350 203008 334384
rect 202688 334294 202758 334350
rect 202814 334294 202882 334350
rect 202938 334294 203008 334350
rect 202688 334226 203008 334294
rect 202688 334170 202758 334226
rect 202814 334170 202882 334226
rect 202938 334170 203008 334226
rect 202688 334102 203008 334170
rect 202688 334046 202758 334102
rect 202814 334046 202882 334102
rect 202938 334046 203008 334102
rect 202688 333978 203008 334046
rect 202688 333922 202758 333978
rect 202814 333922 202882 333978
rect 202938 333922 203008 333978
rect 202688 333888 203008 333922
rect 233408 334350 233728 334384
rect 233408 334294 233478 334350
rect 233534 334294 233602 334350
rect 233658 334294 233728 334350
rect 233408 334226 233728 334294
rect 233408 334170 233478 334226
rect 233534 334170 233602 334226
rect 233658 334170 233728 334226
rect 233408 334102 233728 334170
rect 233408 334046 233478 334102
rect 233534 334046 233602 334102
rect 233658 334046 233728 334102
rect 233408 333978 233728 334046
rect 233408 333922 233478 333978
rect 233534 333922 233602 333978
rect 233658 333922 233728 333978
rect 233408 333888 233728 333922
rect 264128 334350 264448 334384
rect 264128 334294 264198 334350
rect 264254 334294 264322 334350
rect 264378 334294 264448 334350
rect 264128 334226 264448 334294
rect 264128 334170 264198 334226
rect 264254 334170 264322 334226
rect 264378 334170 264448 334226
rect 264128 334102 264448 334170
rect 264128 334046 264198 334102
rect 264254 334046 264322 334102
rect 264378 334046 264448 334102
rect 264128 333978 264448 334046
rect 264128 333922 264198 333978
rect 264254 333922 264322 333978
rect 264378 333922 264448 333978
rect 264128 333888 264448 333922
rect 294848 334350 295168 334384
rect 294848 334294 294918 334350
rect 294974 334294 295042 334350
rect 295098 334294 295168 334350
rect 294848 334226 295168 334294
rect 294848 334170 294918 334226
rect 294974 334170 295042 334226
rect 295098 334170 295168 334226
rect 294848 334102 295168 334170
rect 294848 334046 294918 334102
rect 294974 334046 295042 334102
rect 295098 334046 295168 334102
rect 294848 333978 295168 334046
rect 294848 333922 294918 333978
rect 294974 333922 295042 333978
rect 295098 333922 295168 333978
rect 294848 333888 295168 333922
rect 325568 334350 325888 334384
rect 325568 334294 325638 334350
rect 325694 334294 325762 334350
rect 325818 334294 325888 334350
rect 325568 334226 325888 334294
rect 325568 334170 325638 334226
rect 325694 334170 325762 334226
rect 325818 334170 325888 334226
rect 325568 334102 325888 334170
rect 325568 334046 325638 334102
rect 325694 334046 325762 334102
rect 325818 334046 325888 334102
rect 325568 333978 325888 334046
rect 325568 333922 325638 333978
rect 325694 333922 325762 333978
rect 325818 333922 325888 333978
rect 325568 333888 325888 333922
rect 348874 334350 349494 351922
rect 356288 352350 356608 352384
rect 356288 352294 356358 352350
rect 356414 352294 356482 352350
rect 356538 352294 356608 352350
rect 356288 352226 356608 352294
rect 356288 352170 356358 352226
rect 356414 352170 356482 352226
rect 356538 352170 356608 352226
rect 356288 352102 356608 352170
rect 356288 352046 356358 352102
rect 356414 352046 356482 352102
rect 356538 352046 356608 352102
rect 356288 351978 356608 352046
rect 356288 351922 356358 351978
rect 356414 351922 356482 351978
rect 356538 351922 356608 351978
rect 356288 351888 356608 351922
rect 363154 346350 363774 363922
rect 363154 346294 363250 346350
rect 363306 346294 363374 346350
rect 363430 346294 363498 346350
rect 363554 346294 363622 346350
rect 363678 346294 363774 346350
rect 363154 346226 363774 346294
rect 363154 346170 363250 346226
rect 363306 346170 363374 346226
rect 363430 346170 363498 346226
rect 363554 346170 363622 346226
rect 363678 346170 363774 346226
rect 363154 346102 363774 346170
rect 363154 346046 363250 346102
rect 363306 346046 363374 346102
rect 363430 346046 363498 346102
rect 363554 346046 363622 346102
rect 363678 346046 363774 346102
rect 363154 345978 363774 346046
rect 363154 345922 363250 345978
rect 363306 345922 363374 345978
rect 363430 345922 363498 345978
rect 363554 345922 363622 345978
rect 363678 345922 363774 345978
rect 348874 334294 348970 334350
rect 349026 334294 349094 334350
rect 349150 334294 349218 334350
rect 349274 334294 349342 334350
rect 349398 334294 349494 334350
rect 348874 334226 349494 334294
rect 348874 334170 348970 334226
rect 349026 334170 349094 334226
rect 349150 334170 349218 334226
rect 349274 334170 349342 334226
rect 349398 334170 349494 334226
rect 348874 334102 349494 334170
rect 348874 334046 348970 334102
rect 349026 334046 349094 334102
rect 349150 334046 349218 334102
rect 349274 334046 349342 334102
rect 349398 334046 349494 334102
rect 348874 333978 349494 334046
rect 348874 333922 348970 333978
rect 349026 333922 349094 333978
rect 349150 333922 349218 333978
rect 349274 333922 349342 333978
rect 349398 333922 349494 333978
rect 57154 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 57774 328350
rect 57154 328226 57774 328294
rect 57154 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 57774 328226
rect 57154 328102 57774 328170
rect 57154 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 57774 328102
rect 57154 327978 57774 328046
rect 57154 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 57774 327978
rect 57154 310350 57774 327922
rect 64448 328350 64768 328384
rect 64448 328294 64518 328350
rect 64574 328294 64642 328350
rect 64698 328294 64768 328350
rect 64448 328226 64768 328294
rect 64448 328170 64518 328226
rect 64574 328170 64642 328226
rect 64698 328170 64768 328226
rect 64448 328102 64768 328170
rect 64448 328046 64518 328102
rect 64574 328046 64642 328102
rect 64698 328046 64768 328102
rect 64448 327978 64768 328046
rect 64448 327922 64518 327978
rect 64574 327922 64642 327978
rect 64698 327922 64768 327978
rect 64448 327888 64768 327922
rect 95168 328350 95488 328384
rect 95168 328294 95238 328350
rect 95294 328294 95362 328350
rect 95418 328294 95488 328350
rect 95168 328226 95488 328294
rect 95168 328170 95238 328226
rect 95294 328170 95362 328226
rect 95418 328170 95488 328226
rect 95168 328102 95488 328170
rect 95168 328046 95238 328102
rect 95294 328046 95362 328102
rect 95418 328046 95488 328102
rect 95168 327978 95488 328046
rect 95168 327922 95238 327978
rect 95294 327922 95362 327978
rect 95418 327922 95488 327978
rect 95168 327888 95488 327922
rect 125888 328350 126208 328384
rect 125888 328294 125958 328350
rect 126014 328294 126082 328350
rect 126138 328294 126208 328350
rect 125888 328226 126208 328294
rect 125888 328170 125958 328226
rect 126014 328170 126082 328226
rect 126138 328170 126208 328226
rect 125888 328102 126208 328170
rect 125888 328046 125958 328102
rect 126014 328046 126082 328102
rect 126138 328046 126208 328102
rect 125888 327978 126208 328046
rect 125888 327922 125958 327978
rect 126014 327922 126082 327978
rect 126138 327922 126208 327978
rect 125888 327888 126208 327922
rect 156608 328350 156928 328384
rect 156608 328294 156678 328350
rect 156734 328294 156802 328350
rect 156858 328294 156928 328350
rect 156608 328226 156928 328294
rect 156608 328170 156678 328226
rect 156734 328170 156802 328226
rect 156858 328170 156928 328226
rect 156608 328102 156928 328170
rect 156608 328046 156678 328102
rect 156734 328046 156802 328102
rect 156858 328046 156928 328102
rect 156608 327978 156928 328046
rect 156608 327922 156678 327978
rect 156734 327922 156802 327978
rect 156858 327922 156928 327978
rect 156608 327888 156928 327922
rect 187328 328350 187648 328384
rect 187328 328294 187398 328350
rect 187454 328294 187522 328350
rect 187578 328294 187648 328350
rect 187328 328226 187648 328294
rect 187328 328170 187398 328226
rect 187454 328170 187522 328226
rect 187578 328170 187648 328226
rect 187328 328102 187648 328170
rect 187328 328046 187398 328102
rect 187454 328046 187522 328102
rect 187578 328046 187648 328102
rect 187328 327978 187648 328046
rect 187328 327922 187398 327978
rect 187454 327922 187522 327978
rect 187578 327922 187648 327978
rect 187328 327888 187648 327922
rect 218048 328350 218368 328384
rect 218048 328294 218118 328350
rect 218174 328294 218242 328350
rect 218298 328294 218368 328350
rect 218048 328226 218368 328294
rect 218048 328170 218118 328226
rect 218174 328170 218242 328226
rect 218298 328170 218368 328226
rect 218048 328102 218368 328170
rect 218048 328046 218118 328102
rect 218174 328046 218242 328102
rect 218298 328046 218368 328102
rect 218048 327978 218368 328046
rect 218048 327922 218118 327978
rect 218174 327922 218242 327978
rect 218298 327922 218368 327978
rect 218048 327888 218368 327922
rect 248768 328350 249088 328384
rect 248768 328294 248838 328350
rect 248894 328294 248962 328350
rect 249018 328294 249088 328350
rect 248768 328226 249088 328294
rect 248768 328170 248838 328226
rect 248894 328170 248962 328226
rect 249018 328170 249088 328226
rect 248768 328102 249088 328170
rect 248768 328046 248838 328102
rect 248894 328046 248962 328102
rect 249018 328046 249088 328102
rect 248768 327978 249088 328046
rect 248768 327922 248838 327978
rect 248894 327922 248962 327978
rect 249018 327922 249088 327978
rect 248768 327888 249088 327922
rect 279488 328350 279808 328384
rect 279488 328294 279558 328350
rect 279614 328294 279682 328350
rect 279738 328294 279808 328350
rect 279488 328226 279808 328294
rect 279488 328170 279558 328226
rect 279614 328170 279682 328226
rect 279738 328170 279808 328226
rect 279488 328102 279808 328170
rect 279488 328046 279558 328102
rect 279614 328046 279682 328102
rect 279738 328046 279808 328102
rect 279488 327978 279808 328046
rect 279488 327922 279558 327978
rect 279614 327922 279682 327978
rect 279738 327922 279808 327978
rect 279488 327888 279808 327922
rect 310208 328350 310528 328384
rect 310208 328294 310278 328350
rect 310334 328294 310402 328350
rect 310458 328294 310528 328350
rect 310208 328226 310528 328294
rect 310208 328170 310278 328226
rect 310334 328170 310402 328226
rect 310458 328170 310528 328226
rect 310208 328102 310528 328170
rect 310208 328046 310278 328102
rect 310334 328046 310402 328102
rect 310458 328046 310528 328102
rect 310208 327978 310528 328046
rect 310208 327922 310278 327978
rect 310334 327922 310402 327978
rect 310458 327922 310528 327978
rect 310208 327888 310528 327922
rect 340928 328350 341248 328384
rect 340928 328294 340998 328350
rect 341054 328294 341122 328350
rect 341178 328294 341248 328350
rect 340928 328226 341248 328294
rect 340928 328170 340998 328226
rect 341054 328170 341122 328226
rect 341178 328170 341248 328226
rect 340928 328102 341248 328170
rect 340928 328046 340998 328102
rect 341054 328046 341122 328102
rect 341178 328046 341248 328102
rect 340928 327978 341248 328046
rect 340928 327922 340998 327978
rect 341054 327922 341122 327978
rect 341178 327922 341248 327978
rect 340928 327888 341248 327922
rect 79808 316350 80128 316384
rect 79808 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 80128 316350
rect 79808 316226 80128 316294
rect 79808 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 80128 316226
rect 79808 316102 80128 316170
rect 79808 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 80128 316102
rect 79808 315978 80128 316046
rect 79808 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 80128 315978
rect 79808 315888 80128 315922
rect 110528 316350 110848 316384
rect 110528 316294 110598 316350
rect 110654 316294 110722 316350
rect 110778 316294 110848 316350
rect 110528 316226 110848 316294
rect 110528 316170 110598 316226
rect 110654 316170 110722 316226
rect 110778 316170 110848 316226
rect 110528 316102 110848 316170
rect 110528 316046 110598 316102
rect 110654 316046 110722 316102
rect 110778 316046 110848 316102
rect 110528 315978 110848 316046
rect 110528 315922 110598 315978
rect 110654 315922 110722 315978
rect 110778 315922 110848 315978
rect 110528 315888 110848 315922
rect 141248 316350 141568 316384
rect 141248 316294 141318 316350
rect 141374 316294 141442 316350
rect 141498 316294 141568 316350
rect 141248 316226 141568 316294
rect 141248 316170 141318 316226
rect 141374 316170 141442 316226
rect 141498 316170 141568 316226
rect 141248 316102 141568 316170
rect 141248 316046 141318 316102
rect 141374 316046 141442 316102
rect 141498 316046 141568 316102
rect 141248 315978 141568 316046
rect 141248 315922 141318 315978
rect 141374 315922 141442 315978
rect 141498 315922 141568 315978
rect 141248 315888 141568 315922
rect 171968 316350 172288 316384
rect 171968 316294 172038 316350
rect 172094 316294 172162 316350
rect 172218 316294 172288 316350
rect 171968 316226 172288 316294
rect 171968 316170 172038 316226
rect 172094 316170 172162 316226
rect 172218 316170 172288 316226
rect 171968 316102 172288 316170
rect 171968 316046 172038 316102
rect 172094 316046 172162 316102
rect 172218 316046 172288 316102
rect 171968 315978 172288 316046
rect 171968 315922 172038 315978
rect 172094 315922 172162 315978
rect 172218 315922 172288 315978
rect 171968 315888 172288 315922
rect 202688 316350 203008 316384
rect 202688 316294 202758 316350
rect 202814 316294 202882 316350
rect 202938 316294 203008 316350
rect 202688 316226 203008 316294
rect 202688 316170 202758 316226
rect 202814 316170 202882 316226
rect 202938 316170 203008 316226
rect 202688 316102 203008 316170
rect 202688 316046 202758 316102
rect 202814 316046 202882 316102
rect 202938 316046 203008 316102
rect 202688 315978 203008 316046
rect 202688 315922 202758 315978
rect 202814 315922 202882 315978
rect 202938 315922 203008 315978
rect 202688 315888 203008 315922
rect 233408 316350 233728 316384
rect 233408 316294 233478 316350
rect 233534 316294 233602 316350
rect 233658 316294 233728 316350
rect 233408 316226 233728 316294
rect 233408 316170 233478 316226
rect 233534 316170 233602 316226
rect 233658 316170 233728 316226
rect 233408 316102 233728 316170
rect 233408 316046 233478 316102
rect 233534 316046 233602 316102
rect 233658 316046 233728 316102
rect 233408 315978 233728 316046
rect 233408 315922 233478 315978
rect 233534 315922 233602 315978
rect 233658 315922 233728 315978
rect 233408 315888 233728 315922
rect 264128 316350 264448 316384
rect 264128 316294 264198 316350
rect 264254 316294 264322 316350
rect 264378 316294 264448 316350
rect 264128 316226 264448 316294
rect 264128 316170 264198 316226
rect 264254 316170 264322 316226
rect 264378 316170 264448 316226
rect 264128 316102 264448 316170
rect 264128 316046 264198 316102
rect 264254 316046 264322 316102
rect 264378 316046 264448 316102
rect 264128 315978 264448 316046
rect 264128 315922 264198 315978
rect 264254 315922 264322 315978
rect 264378 315922 264448 315978
rect 264128 315888 264448 315922
rect 294848 316350 295168 316384
rect 294848 316294 294918 316350
rect 294974 316294 295042 316350
rect 295098 316294 295168 316350
rect 294848 316226 295168 316294
rect 294848 316170 294918 316226
rect 294974 316170 295042 316226
rect 295098 316170 295168 316226
rect 294848 316102 295168 316170
rect 294848 316046 294918 316102
rect 294974 316046 295042 316102
rect 295098 316046 295168 316102
rect 294848 315978 295168 316046
rect 294848 315922 294918 315978
rect 294974 315922 295042 315978
rect 295098 315922 295168 315978
rect 294848 315888 295168 315922
rect 325568 316350 325888 316384
rect 325568 316294 325638 316350
rect 325694 316294 325762 316350
rect 325818 316294 325888 316350
rect 325568 316226 325888 316294
rect 325568 316170 325638 316226
rect 325694 316170 325762 316226
rect 325818 316170 325888 316226
rect 325568 316102 325888 316170
rect 325568 316046 325638 316102
rect 325694 316046 325762 316102
rect 325818 316046 325888 316102
rect 325568 315978 325888 316046
rect 325568 315922 325638 315978
rect 325694 315922 325762 315978
rect 325818 315922 325888 315978
rect 325568 315888 325888 315922
rect 348874 316350 349494 333922
rect 356288 334350 356608 334384
rect 356288 334294 356358 334350
rect 356414 334294 356482 334350
rect 356538 334294 356608 334350
rect 356288 334226 356608 334294
rect 356288 334170 356358 334226
rect 356414 334170 356482 334226
rect 356538 334170 356608 334226
rect 356288 334102 356608 334170
rect 356288 334046 356358 334102
rect 356414 334046 356482 334102
rect 356538 334046 356608 334102
rect 356288 333978 356608 334046
rect 356288 333922 356358 333978
rect 356414 333922 356482 333978
rect 356538 333922 356608 333978
rect 356288 333888 356608 333922
rect 363154 328350 363774 345922
rect 363154 328294 363250 328350
rect 363306 328294 363374 328350
rect 363430 328294 363498 328350
rect 363554 328294 363622 328350
rect 363678 328294 363774 328350
rect 363154 328226 363774 328294
rect 363154 328170 363250 328226
rect 363306 328170 363374 328226
rect 363430 328170 363498 328226
rect 363554 328170 363622 328226
rect 363678 328170 363774 328226
rect 363154 328102 363774 328170
rect 363154 328046 363250 328102
rect 363306 328046 363374 328102
rect 363430 328046 363498 328102
rect 363554 328046 363622 328102
rect 363678 328046 363774 328102
rect 363154 327978 363774 328046
rect 363154 327922 363250 327978
rect 363306 327922 363374 327978
rect 363430 327922 363498 327978
rect 363554 327922 363622 327978
rect 363678 327922 363774 327978
rect 348874 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 349494 316350
rect 348874 316226 349494 316294
rect 348874 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 349494 316226
rect 348874 316102 349494 316170
rect 348874 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 349494 316102
rect 348874 315978 349494 316046
rect 348874 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 349494 315978
rect 57154 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 57774 310350
rect 57154 310226 57774 310294
rect 57154 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 57774 310226
rect 57154 310102 57774 310170
rect 57154 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 57774 310102
rect 57154 309978 57774 310046
rect 57154 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 57774 309978
rect 57154 292350 57774 309922
rect 64448 310350 64768 310384
rect 64448 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 64768 310350
rect 64448 310226 64768 310294
rect 64448 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 64768 310226
rect 64448 310102 64768 310170
rect 64448 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 64768 310102
rect 64448 309978 64768 310046
rect 64448 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 64768 309978
rect 64448 309888 64768 309922
rect 95168 310350 95488 310384
rect 95168 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 95488 310350
rect 95168 310226 95488 310294
rect 95168 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 95488 310226
rect 95168 310102 95488 310170
rect 95168 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 95488 310102
rect 95168 309978 95488 310046
rect 95168 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 95488 309978
rect 95168 309888 95488 309922
rect 125888 310350 126208 310384
rect 125888 310294 125958 310350
rect 126014 310294 126082 310350
rect 126138 310294 126208 310350
rect 125888 310226 126208 310294
rect 125888 310170 125958 310226
rect 126014 310170 126082 310226
rect 126138 310170 126208 310226
rect 125888 310102 126208 310170
rect 125888 310046 125958 310102
rect 126014 310046 126082 310102
rect 126138 310046 126208 310102
rect 125888 309978 126208 310046
rect 125888 309922 125958 309978
rect 126014 309922 126082 309978
rect 126138 309922 126208 309978
rect 125888 309888 126208 309922
rect 156608 310350 156928 310384
rect 156608 310294 156678 310350
rect 156734 310294 156802 310350
rect 156858 310294 156928 310350
rect 156608 310226 156928 310294
rect 156608 310170 156678 310226
rect 156734 310170 156802 310226
rect 156858 310170 156928 310226
rect 156608 310102 156928 310170
rect 156608 310046 156678 310102
rect 156734 310046 156802 310102
rect 156858 310046 156928 310102
rect 156608 309978 156928 310046
rect 156608 309922 156678 309978
rect 156734 309922 156802 309978
rect 156858 309922 156928 309978
rect 156608 309888 156928 309922
rect 187328 310350 187648 310384
rect 187328 310294 187398 310350
rect 187454 310294 187522 310350
rect 187578 310294 187648 310350
rect 187328 310226 187648 310294
rect 187328 310170 187398 310226
rect 187454 310170 187522 310226
rect 187578 310170 187648 310226
rect 187328 310102 187648 310170
rect 187328 310046 187398 310102
rect 187454 310046 187522 310102
rect 187578 310046 187648 310102
rect 187328 309978 187648 310046
rect 187328 309922 187398 309978
rect 187454 309922 187522 309978
rect 187578 309922 187648 309978
rect 187328 309888 187648 309922
rect 218048 310350 218368 310384
rect 218048 310294 218118 310350
rect 218174 310294 218242 310350
rect 218298 310294 218368 310350
rect 218048 310226 218368 310294
rect 218048 310170 218118 310226
rect 218174 310170 218242 310226
rect 218298 310170 218368 310226
rect 218048 310102 218368 310170
rect 218048 310046 218118 310102
rect 218174 310046 218242 310102
rect 218298 310046 218368 310102
rect 218048 309978 218368 310046
rect 218048 309922 218118 309978
rect 218174 309922 218242 309978
rect 218298 309922 218368 309978
rect 218048 309888 218368 309922
rect 248768 310350 249088 310384
rect 248768 310294 248838 310350
rect 248894 310294 248962 310350
rect 249018 310294 249088 310350
rect 248768 310226 249088 310294
rect 248768 310170 248838 310226
rect 248894 310170 248962 310226
rect 249018 310170 249088 310226
rect 248768 310102 249088 310170
rect 248768 310046 248838 310102
rect 248894 310046 248962 310102
rect 249018 310046 249088 310102
rect 248768 309978 249088 310046
rect 248768 309922 248838 309978
rect 248894 309922 248962 309978
rect 249018 309922 249088 309978
rect 248768 309888 249088 309922
rect 279488 310350 279808 310384
rect 279488 310294 279558 310350
rect 279614 310294 279682 310350
rect 279738 310294 279808 310350
rect 279488 310226 279808 310294
rect 279488 310170 279558 310226
rect 279614 310170 279682 310226
rect 279738 310170 279808 310226
rect 279488 310102 279808 310170
rect 279488 310046 279558 310102
rect 279614 310046 279682 310102
rect 279738 310046 279808 310102
rect 279488 309978 279808 310046
rect 279488 309922 279558 309978
rect 279614 309922 279682 309978
rect 279738 309922 279808 309978
rect 279488 309888 279808 309922
rect 310208 310350 310528 310384
rect 310208 310294 310278 310350
rect 310334 310294 310402 310350
rect 310458 310294 310528 310350
rect 310208 310226 310528 310294
rect 310208 310170 310278 310226
rect 310334 310170 310402 310226
rect 310458 310170 310528 310226
rect 310208 310102 310528 310170
rect 310208 310046 310278 310102
rect 310334 310046 310402 310102
rect 310458 310046 310528 310102
rect 310208 309978 310528 310046
rect 310208 309922 310278 309978
rect 310334 309922 310402 309978
rect 310458 309922 310528 309978
rect 310208 309888 310528 309922
rect 340928 310350 341248 310384
rect 340928 310294 340998 310350
rect 341054 310294 341122 310350
rect 341178 310294 341248 310350
rect 340928 310226 341248 310294
rect 340928 310170 340998 310226
rect 341054 310170 341122 310226
rect 341178 310170 341248 310226
rect 340928 310102 341248 310170
rect 340928 310046 340998 310102
rect 341054 310046 341122 310102
rect 341178 310046 341248 310102
rect 340928 309978 341248 310046
rect 340928 309922 340998 309978
rect 341054 309922 341122 309978
rect 341178 309922 341248 309978
rect 340928 309888 341248 309922
rect 79808 298350 80128 298384
rect 79808 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 80128 298350
rect 79808 298226 80128 298294
rect 79808 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 80128 298226
rect 79808 298102 80128 298170
rect 79808 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 80128 298102
rect 79808 297978 80128 298046
rect 79808 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 80128 297978
rect 79808 297888 80128 297922
rect 110528 298350 110848 298384
rect 110528 298294 110598 298350
rect 110654 298294 110722 298350
rect 110778 298294 110848 298350
rect 110528 298226 110848 298294
rect 110528 298170 110598 298226
rect 110654 298170 110722 298226
rect 110778 298170 110848 298226
rect 110528 298102 110848 298170
rect 110528 298046 110598 298102
rect 110654 298046 110722 298102
rect 110778 298046 110848 298102
rect 110528 297978 110848 298046
rect 110528 297922 110598 297978
rect 110654 297922 110722 297978
rect 110778 297922 110848 297978
rect 110528 297888 110848 297922
rect 141248 298350 141568 298384
rect 141248 298294 141318 298350
rect 141374 298294 141442 298350
rect 141498 298294 141568 298350
rect 141248 298226 141568 298294
rect 141248 298170 141318 298226
rect 141374 298170 141442 298226
rect 141498 298170 141568 298226
rect 141248 298102 141568 298170
rect 141248 298046 141318 298102
rect 141374 298046 141442 298102
rect 141498 298046 141568 298102
rect 141248 297978 141568 298046
rect 141248 297922 141318 297978
rect 141374 297922 141442 297978
rect 141498 297922 141568 297978
rect 141248 297888 141568 297922
rect 171968 298350 172288 298384
rect 171968 298294 172038 298350
rect 172094 298294 172162 298350
rect 172218 298294 172288 298350
rect 171968 298226 172288 298294
rect 171968 298170 172038 298226
rect 172094 298170 172162 298226
rect 172218 298170 172288 298226
rect 171968 298102 172288 298170
rect 171968 298046 172038 298102
rect 172094 298046 172162 298102
rect 172218 298046 172288 298102
rect 171968 297978 172288 298046
rect 171968 297922 172038 297978
rect 172094 297922 172162 297978
rect 172218 297922 172288 297978
rect 171968 297888 172288 297922
rect 202688 298350 203008 298384
rect 202688 298294 202758 298350
rect 202814 298294 202882 298350
rect 202938 298294 203008 298350
rect 202688 298226 203008 298294
rect 202688 298170 202758 298226
rect 202814 298170 202882 298226
rect 202938 298170 203008 298226
rect 202688 298102 203008 298170
rect 202688 298046 202758 298102
rect 202814 298046 202882 298102
rect 202938 298046 203008 298102
rect 202688 297978 203008 298046
rect 202688 297922 202758 297978
rect 202814 297922 202882 297978
rect 202938 297922 203008 297978
rect 202688 297888 203008 297922
rect 233408 298350 233728 298384
rect 233408 298294 233478 298350
rect 233534 298294 233602 298350
rect 233658 298294 233728 298350
rect 233408 298226 233728 298294
rect 233408 298170 233478 298226
rect 233534 298170 233602 298226
rect 233658 298170 233728 298226
rect 233408 298102 233728 298170
rect 233408 298046 233478 298102
rect 233534 298046 233602 298102
rect 233658 298046 233728 298102
rect 233408 297978 233728 298046
rect 233408 297922 233478 297978
rect 233534 297922 233602 297978
rect 233658 297922 233728 297978
rect 233408 297888 233728 297922
rect 264128 298350 264448 298384
rect 264128 298294 264198 298350
rect 264254 298294 264322 298350
rect 264378 298294 264448 298350
rect 264128 298226 264448 298294
rect 264128 298170 264198 298226
rect 264254 298170 264322 298226
rect 264378 298170 264448 298226
rect 264128 298102 264448 298170
rect 264128 298046 264198 298102
rect 264254 298046 264322 298102
rect 264378 298046 264448 298102
rect 264128 297978 264448 298046
rect 264128 297922 264198 297978
rect 264254 297922 264322 297978
rect 264378 297922 264448 297978
rect 264128 297888 264448 297922
rect 294848 298350 295168 298384
rect 294848 298294 294918 298350
rect 294974 298294 295042 298350
rect 295098 298294 295168 298350
rect 294848 298226 295168 298294
rect 294848 298170 294918 298226
rect 294974 298170 295042 298226
rect 295098 298170 295168 298226
rect 294848 298102 295168 298170
rect 294848 298046 294918 298102
rect 294974 298046 295042 298102
rect 295098 298046 295168 298102
rect 294848 297978 295168 298046
rect 294848 297922 294918 297978
rect 294974 297922 295042 297978
rect 295098 297922 295168 297978
rect 294848 297888 295168 297922
rect 325568 298350 325888 298384
rect 325568 298294 325638 298350
rect 325694 298294 325762 298350
rect 325818 298294 325888 298350
rect 325568 298226 325888 298294
rect 325568 298170 325638 298226
rect 325694 298170 325762 298226
rect 325818 298170 325888 298226
rect 325568 298102 325888 298170
rect 325568 298046 325638 298102
rect 325694 298046 325762 298102
rect 325818 298046 325888 298102
rect 325568 297978 325888 298046
rect 325568 297922 325638 297978
rect 325694 297922 325762 297978
rect 325818 297922 325888 297978
rect 325568 297888 325888 297922
rect 348874 298350 349494 315922
rect 356288 316350 356608 316384
rect 356288 316294 356358 316350
rect 356414 316294 356482 316350
rect 356538 316294 356608 316350
rect 356288 316226 356608 316294
rect 356288 316170 356358 316226
rect 356414 316170 356482 316226
rect 356538 316170 356608 316226
rect 356288 316102 356608 316170
rect 356288 316046 356358 316102
rect 356414 316046 356482 316102
rect 356538 316046 356608 316102
rect 356288 315978 356608 316046
rect 356288 315922 356358 315978
rect 356414 315922 356482 315978
rect 356538 315922 356608 315978
rect 356288 315888 356608 315922
rect 363154 310350 363774 327922
rect 363154 310294 363250 310350
rect 363306 310294 363374 310350
rect 363430 310294 363498 310350
rect 363554 310294 363622 310350
rect 363678 310294 363774 310350
rect 363154 310226 363774 310294
rect 363154 310170 363250 310226
rect 363306 310170 363374 310226
rect 363430 310170 363498 310226
rect 363554 310170 363622 310226
rect 363678 310170 363774 310226
rect 363154 310102 363774 310170
rect 363154 310046 363250 310102
rect 363306 310046 363374 310102
rect 363430 310046 363498 310102
rect 363554 310046 363622 310102
rect 363678 310046 363774 310102
rect 363154 309978 363774 310046
rect 363154 309922 363250 309978
rect 363306 309922 363374 309978
rect 363430 309922 363498 309978
rect 363554 309922 363622 309978
rect 363678 309922 363774 309978
rect 348874 298294 348970 298350
rect 349026 298294 349094 298350
rect 349150 298294 349218 298350
rect 349274 298294 349342 298350
rect 349398 298294 349494 298350
rect 348874 298226 349494 298294
rect 348874 298170 348970 298226
rect 349026 298170 349094 298226
rect 349150 298170 349218 298226
rect 349274 298170 349342 298226
rect 349398 298170 349494 298226
rect 348874 298102 349494 298170
rect 348874 298046 348970 298102
rect 349026 298046 349094 298102
rect 349150 298046 349218 298102
rect 349274 298046 349342 298102
rect 349398 298046 349494 298102
rect 348874 297978 349494 298046
rect 348874 297922 348970 297978
rect 349026 297922 349094 297978
rect 349150 297922 349218 297978
rect 349274 297922 349342 297978
rect 349398 297922 349494 297978
rect 57154 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 57774 292350
rect 57154 292226 57774 292294
rect 57154 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 57774 292226
rect 57154 292102 57774 292170
rect 57154 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 57774 292102
rect 57154 291978 57774 292046
rect 57154 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 57774 291978
rect 57154 274350 57774 291922
rect 64448 292350 64768 292384
rect 64448 292294 64518 292350
rect 64574 292294 64642 292350
rect 64698 292294 64768 292350
rect 64448 292226 64768 292294
rect 64448 292170 64518 292226
rect 64574 292170 64642 292226
rect 64698 292170 64768 292226
rect 64448 292102 64768 292170
rect 64448 292046 64518 292102
rect 64574 292046 64642 292102
rect 64698 292046 64768 292102
rect 64448 291978 64768 292046
rect 64448 291922 64518 291978
rect 64574 291922 64642 291978
rect 64698 291922 64768 291978
rect 64448 291888 64768 291922
rect 95168 292350 95488 292384
rect 95168 292294 95238 292350
rect 95294 292294 95362 292350
rect 95418 292294 95488 292350
rect 95168 292226 95488 292294
rect 95168 292170 95238 292226
rect 95294 292170 95362 292226
rect 95418 292170 95488 292226
rect 95168 292102 95488 292170
rect 95168 292046 95238 292102
rect 95294 292046 95362 292102
rect 95418 292046 95488 292102
rect 95168 291978 95488 292046
rect 95168 291922 95238 291978
rect 95294 291922 95362 291978
rect 95418 291922 95488 291978
rect 95168 291888 95488 291922
rect 125888 292350 126208 292384
rect 125888 292294 125958 292350
rect 126014 292294 126082 292350
rect 126138 292294 126208 292350
rect 125888 292226 126208 292294
rect 125888 292170 125958 292226
rect 126014 292170 126082 292226
rect 126138 292170 126208 292226
rect 125888 292102 126208 292170
rect 125888 292046 125958 292102
rect 126014 292046 126082 292102
rect 126138 292046 126208 292102
rect 125888 291978 126208 292046
rect 125888 291922 125958 291978
rect 126014 291922 126082 291978
rect 126138 291922 126208 291978
rect 125888 291888 126208 291922
rect 156608 292350 156928 292384
rect 156608 292294 156678 292350
rect 156734 292294 156802 292350
rect 156858 292294 156928 292350
rect 156608 292226 156928 292294
rect 156608 292170 156678 292226
rect 156734 292170 156802 292226
rect 156858 292170 156928 292226
rect 156608 292102 156928 292170
rect 156608 292046 156678 292102
rect 156734 292046 156802 292102
rect 156858 292046 156928 292102
rect 156608 291978 156928 292046
rect 156608 291922 156678 291978
rect 156734 291922 156802 291978
rect 156858 291922 156928 291978
rect 156608 291888 156928 291922
rect 187328 292350 187648 292384
rect 187328 292294 187398 292350
rect 187454 292294 187522 292350
rect 187578 292294 187648 292350
rect 187328 292226 187648 292294
rect 187328 292170 187398 292226
rect 187454 292170 187522 292226
rect 187578 292170 187648 292226
rect 187328 292102 187648 292170
rect 187328 292046 187398 292102
rect 187454 292046 187522 292102
rect 187578 292046 187648 292102
rect 187328 291978 187648 292046
rect 187328 291922 187398 291978
rect 187454 291922 187522 291978
rect 187578 291922 187648 291978
rect 187328 291888 187648 291922
rect 218048 292350 218368 292384
rect 218048 292294 218118 292350
rect 218174 292294 218242 292350
rect 218298 292294 218368 292350
rect 218048 292226 218368 292294
rect 218048 292170 218118 292226
rect 218174 292170 218242 292226
rect 218298 292170 218368 292226
rect 218048 292102 218368 292170
rect 218048 292046 218118 292102
rect 218174 292046 218242 292102
rect 218298 292046 218368 292102
rect 218048 291978 218368 292046
rect 218048 291922 218118 291978
rect 218174 291922 218242 291978
rect 218298 291922 218368 291978
rect 218048 291888 218368 291922
rect 248768 292350 249088 292384
rect 248768 292294 248838 292350
rect 248894 292294 248962 292350
rect 249018 292294 249088 292350
rect 248768 292226 249088 292294
rect 248768 292170 248838 292226
rect 248894 292170 248962 292226
rect 249018 292170 249088 292226
rect 248768 292102 249088 292170
rect 248768 292046 248838 292102
rect 248894 292046 248962 292102
rect 249018 292046 249088 292102
rect 248768 291978 249088 292046
rect 248768 291922 248838 291978
rect 248894 291922 248962 291978
rect 249018 291922 249088 291978
rect 248768 291888 249088 291922
rect 279488 292350 279808 292384
rect 279488 292294 279558 292350
rect 279614 292294 279682 292350
rect 279738 292294 279808 292350
rect 279488 292226 279808 292294
rect 279488 292170 279558 292226
rect 279614 292170 279682 292226
rect 279738 292170 279808 292226
rect 279488 292102 279808 292170
rect 279488 292046 279558 292102
rect 279614 292046 279682 292102
rect 279738 292046 279808 292102
rect 279488 291978 279808 292046
rect 279488 291922 279558 291978
rect 279614 291922 279682 291978
rect 279738 291922 279808 291978
rect 279488 291888 279808 291922
rect 310208 292350 310528 292384
rect 310208 292294 310278 292350
rect 310334 292294 310402 292350
rect 310458 292294 310528 292350
rect 310208 292226 310528 292294
rect 310208 292170 310278 292226
rect 310334 292170 310402 292226
rect 310458 292170 310528 292226
rect 310208 292102 310528 292170
rect 310208 292046 310278 292102
rect 310334 292046 310402 292102
rect 310458 292046 310528 292102
rect 310208 291978 310528 292046
rect 310208 291922 310278 291978
rect 310334 291922 310402 291978
rect 310458 291922 310528 291978
rect 310208 291888 310528 291922
rect 340928 292350 341248 292384
rect 340928 292294 340998 292350
rect 341054 292294 341122 292350
rect 341178 292294 341248 292350
rect 340928 292226 341248 292294
rect 340928 292170 340998 292226
rect 341054 292170 341122 292226
rect 341178 292170 341248 292226
rect 340928 292102 341248 292170
rect 340928 292046 340998 292102
rect 341054 292046 341122 292102
rect 341178 292046 341248 292102
rect 340928 291978 341248 292046
rect 340928 291922 340998 291978
rect 341054 291922 341122 291978
rect 341178 291922 341248 291978
rect 340928 291888 341248 291922
rect 79808 280350 80128 280384
rect 79808 280294 79878 280350
rect 79934 280294 80002 280350
rect 80058 280294 80128 280350
rect 79808 280226 80128 280294
rect 79808 280170 79878 280226
rect 79934 280170 80002 280226
rect 80058 280170 80128 280226
rect 79808 280102 80128 280170
rect 79808 280046 79878 280102
rect 79934 280046 80002 280102
rect 80058 280046 80128 280102
rect 79808 279978 80128 280046
rect 79808 279922 79878 279978
rect 79934 279922 80002 279978
rect 80058 279922 80128 279978
rect 79808 279888 80128 279922
rect 110528 280350 110848 280384
rect 110528 280294 110598 280350
rect 110654 280294 110722 280350
rect 110778 280294 110848 280350
rect 110528 280226 110848 280294
rect 110528 280170 110598 280226
rect 110654 280170 110722 280226
rect 110778 280170 110848 280226
rect 110528 280102 110848 280170
rect 110528 280046 110598 280102
rect 110654 280046 110722 280102
rect 110778 280046 110848 280102
rect 110528 279978 110848 280046
rect 110528 279922 110598 279978
rect 110654 279922 110722 279978
rect 110778 279922 110848 279978
rect 110528 279888 110848 279922
rect 141248 280350 141568 280384
rect 141248 280294 141318 280350
rect 141374 280294 141442 280350
rect 141498 280294 141568 280350
rect 141248 280226 141568 280294
rect 141248 280170 141318 280226
rect 141374 280170 141442 280226
rect 141498 280170 141568 280226
rect 141248 280102 141568 280170
rect 141248 280046 141318 280102
rect 141374 280046 141442 280102
rect 141498 280046 141568 280102
rect 141248 279978 141568 280046
rect 141248 279922 141318 279978
rect 141374 279922 141442 279978
rect 141498 279922 141568 279978
rect 141248 279888 141568 279922
rect 171968 280350 172288 280384
rect 171968 280294 172038 280350
rect 172094 280294 172162 280350
rect 172218 280294 172288 280350
rect 171968 280226 172288 280294
rect 171968 280170 172038 280226
rect 172094 280170 172162 280226
rect 172218 280170 172288 280226
rect 171968 280102 172288 280170
rect 171968 280046 172038 280102
rect 172094 280046 172162 280102
rect 172218 280046 172288 280102
rect 171968 279978 172288 280046
rect 171968 279922 172038 279978
rect 172094 279922 172162 279978
rect 172218 279922 172288 279978
rect 171968 279888 172288 279922
rect 202688 280350 203008 280384
rect 202688 280294 202758 280350
rect 202814 280294 202882 280350
rect 202938 280294 203008 280350
rect 202688 280226 203008 280294
rect 202688 280170 202758 280226
rect 202814 280170 202882 280226
rect 202938 280170 203008 280226
rect 202688 280102 203008 280170
rect 202688 280046 202758 280102
rect 202814 280046 202882 280102
rect 202938 280046 203008 280102
rect 202688 279978 203008 280046
rect 202688 279922 202758 279978
rect 202814 279922 202882 279978
rect 202938 279922 203008 279978
rect 202688 279888 203008 279922
rect 233408 280350 233728 280384
rect 233408 280294 233478 280350
rect 233534 280294 233602 280350
rect 233658 280294 233728 280350
rect 233408 280226 233728 280294
rect 233408 280170 233478 280226
rect 233534 280170 233602 280226
rect 233658 280170 233728 280226
rect 233408 280102 233728 280170
rect 233408 280046 233478 280102
rect 233534 280046 233602 280102
rect 233658 280046 233728 280102
rect 233408 279978 233728 280046
rect 233408 279922 233478 279978
rect 233534 279922 233602 279978
rect 233658 279922 233728 279978
rect 233408 279888 233728 279922
rect 264128 280350 264448 280384
rect 264128 280294 264198 280350
rect 264254 280294 264322 280350
rect 264378 280294 264448 280350
rect 264128 280226 264448 280294
rect 264128 280170 264198 280226
rect 264254 280170 264322 280226
rect 264378 280170 264448 280226
rect 264128 280102 264448 280170
rect 264128 280046 264198 280102
rect 264254 280046 264322 280102
rect 264378 280046 264448 280102
rect 264128 279978 264448 280046
rect 264128 279922 264198 279978
rect 264254 279922 264322 279978
rect 264378 279922 264448 279978
rect 264128 279888 264448 279922
rect 294848 280350 295168 280384
rect 294848 280294 294918 280350
rect 294974 280294 295042 280350
rect 295098 280294 295168 280350
rect 294848 280226 295168 280294
rect 294848 280170 294918 280226
rect 294974 280170 295042 280226
rect 295098 280170 295168 280226
rect 294848 280102 295168 280170
rect 294848 280046 294918 280102
rect 294974 280046 295042 280102
rect 295098 280046 295168 280102
rect 294848 279978 295168 280046
rect 294848 279922 294918 279978
rect 294974 279922 295042 279978
rect 295098 279922 295168 279978
rect 294848 279888 295168 279922
rect 325568 280350 325888 280384
rect 325568 280294 325638 280350
rect 325694 280294 325762 280350
rect 325818 280294 325888 280350
rect 325568 280226 325888 280294
rect 325568 280170 325638 280226
rect 325694 280170 325762 280226
rect 325818 280170 325888 280226
rect 325568 280102 325888 280170
rect 325568 280046 325638 280102
rect 325694 280046 325762 280102
rect 325818 280046 325888 280102
rect 325568 279978 325888 280046
rect 325568 279922 325638 279978
rect 325694 279922 325762 279978
rect 325818 279922 325888 279978
rect 325568 279888 325888 279922
rect 348874 280350 349494 297922
rect 356288 298350 356608 298384
rect 356288 298294 356358 298350
rect 356414 298294 356482 298350
rect 356538 298294 356608 298350
rect 356288 298226 356608 298294
rect 356288 298170 356358 298226
rect 356414 298170 356482 298226
rect 356538 298170 356608 298226
rect 356288 298102 356608 298170
rect 356288 298046 356358 298102
rect 356414 298046 356482 298102
rect 356538 298046 356608 298102
rect 356288 297978 356608 298046
rect 356288 297922 356358 297978
rect 356414 297922 356482 297978
rect 356538 297922 356608 297978
rect 356288 297888 356608 297922
rect 363154 292350 363774 309922
rect 363154 292294 363250 292350
rect 363306 292294 363374 292350
rect 363430 292294 363498 292350
rect 363554 292294 363622 292350
rect 363678 292294 363774 292350
rect 363154 292226 363774 292294
rect 363154 292170 363250 292226
rect 363306 292170 363374 292226
rect 363430 292170 363498 292226
rect 363554 292170 363622 292226
rect 363678 292170 363774 292226
rect 363154 292102 363774 292170
rect 363154 292046 363250 292102
rect 363306 292046 363374 292102
rect 363430 292046 363498 292102
rect 363554 292046 363622 292102
rect 363678 292046 363774 292102
rect 363154 291978 363774 292046
rect 363154 291922 363250 291978
rect 363306 291922 363374 291978
rect 363430 291922 363498 291978
rect 363554 291922 363622 291978
rect 363678 291922 363774 291978
rect 348874 280294 348970 280350
rect 349026 280294 349094 280350
rect 349150 280294 349218 280350
rect 349274 280294 349342 280350
rect 349398 280294 349494 280350
rect 348874 280226 349494 280294
rect 348874 280170 348970 280226
rect 349026 280170 349094 280226
rect 349150 280170 349218 280226
rect 349274 280170 349342 280226
rect 349398 280170 349494 280226
rect 348874 280102 349494 280170
rect 348874 280046 348970 280102
rect 349026 280046 349094 280102
rect 349150 280046 349218 280102
rect 349274 280046 349342 280102
rect 349398 280046 349494 280102
rect 348874 279978 349494 280046
rect 348874 279922 348970 279978
rect 349026 279922 349094 279978
rect 349150 279922 349218 279978
rect 349274 279922 349342 279978
rect 349398 279922 349494 279978
rect 57154 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 57774 274350
rect 57154 274226 57774 274294
rect 57154 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 57774 274226
rect 57154 274102 57774 274170
rect 57154 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 57774 274102
rect 57154 273978 57774 274046
rect 57154 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 57774 273978
rect 57154 256350 57774 273922
rect 64448 274350 64768 274384
rect 64448 274294 64518 274350
rect 64574 274294 64642 274350
rect 64698 274294 64768 274350
rect 64448 274226 64768 274294
rect 64448 274170 64518 274226
rect 64574 274170 64642 274226
rect 64698 274170 64768 274226
rect 64448 274102 64768 274170
rect 64448 274046 64518 274102
rect 64574 274046 64642 274102
rect 64698 274046 64768 274102
rect 64448 273978 64768 274046
rect 64448 273922 64518 273978
rect 64574 273922 64642 273978
rect 64698 273922 64768 273978
rect 64448 273888 64768 273922
rect 95168 274350 95488 274384
rect 95168 274294 95238 274350
rect 95294 274294 95362 274350
rect 95418 274294 95488 274350
rect 95168 274226 95488 274294
rect 95168 274170 95238 274226
rect 95294 274170 95362 274226
rect 95418 274170 95488 274226
rect 95168 274102 95488 274170
rect 95168 274046 95238 274102
rect 95294 274046 95362 274102
rect 95418 274046 95488 274102
rect 95168 273978 95488 274046
rect 95168 273922 95238 273978
rect 95294 273922 95362 273978
rect 95418 273922 95488 273978
rect 95168 273888 95488 273922
rect 125888 274350 126208 274384
rect 125888 274294 125958 274350
rect 126014 274294 126082 274350
rect 126138 274294 126208 274350
rect 125888 274226 126208 274294
rect 125888 274170 125958 274226
rect 126014 274170 126082 274226
rect 126138 274170 126208 274226
rect 125888 274102 126208 274170
rect 125888 274046 125958 274102
rect 126014 274046 126082 274102
rect 126138 274046 126208 274102
rect 125888 273978 126208 274046
rect 125888 273922 125958 273978
rect 126014 273922 126082 273978
rect 126138 273922 126208 273978
rect 125888 273888 126208 273922
rect 156608 274350 156928 274384
rect 156608 274294 156678 274350
rect 156734 274294 156802 274350
rect 156858 274294 156928 274350
rect 156608 274226 156928 274294
rect 156608 274170 156678 274226
rect 156734 274170 156802 274226
rect 156858 274170 156928 274226
rect 156608 274102 156928 274170
rect 156608 274046 156678 274102
rect 156734 274046 156802 274102
rect 156858 274046 156928 274102
rect 156608 273978 156928 274046
rect 156608 273922 156678 273978
rect 156734 273922 156802 273978
rect 156858 273922 156928 273978
rect 156608 273888 156928 273922
rect 187328 274350 187648 274384
rect 187328 274294 187398 274350
rect 187454 274294 187522 274350
rect 187578 274294 187648 274350
rect 187328 274226 187648 274294
rect 187328 274170 187398 274226
rect 187454 274170 187522 274226
rect 187578 274170 187648 274226
rect 187328 274102 187648 274170
rect 187328 274046 187398 274102
rect 187454 274046 187522 274102
rect 187578 274046 187648 274102
rect 187328 273978 187648 274046
rect 187328 273922 187398 273978
rect 187454 273922 187522 273978
rect 187578 273922 187648 273978
rect 187328 273888 187648 273922
rect 218048 274350 218368 274384
rect 218048 274294 218118 274350
rect 218174 274294 218242 274350
rect 218298 274294 218368 274350
rect 218048 274226 218368 274294
rect 218048 274170 218118 274226
rect 218174 274170 218242 274226
rect 218298 274170 218368 274226
rect 218048 274102 218368 274170
rect 218048 274046 218118 274102
rect 218174 274046 218242 274102
rect 218298 274046 218368 274102
rect 218048 273978 218368 274046
rect 218048 273922 218118 273978
rect 218174 273922 218242 273978
rect 218298 273922 218368 273978
rect 218048 273888 218368 273922
rect 248768 274350 249088 274384
rect 248768 274294 248838 274350
rect 248894 274294 248962 274350
rect 249018 274294 249088 274350
rect 248768 274226 249088 274294
rect 248768 274170 248838 274226
rect 248894 274170 248962 274226
rect 249018 274170 249088 274226
rect 248768 274102 249088 274170
rect 248768 274046 248838 274102
rect 248894 274046 248962 274102
rect 249018 274046 249088 274102
rect 248768 273978 249088 274046
rect 248768 273922 248838 273978
rect 248894 273922 248962 273978
rect 249018 273922 249088 273978
rect 248768 273888 249088 273922
rect 279488 274350 279808 274384
rect 279488 274294 279558 274350
rect 279614 274294 279682 274350
rect 279738 274294 279808 274350
rect 279488 274226 279808 274294
rect 279488 274170 279558 274226
rect 279614 274170 279682 274226
rect 279738 274170 279808 274226
rect 279488 274102 279808 274170
rect 279488 274046 279558 274102
rect 279614 274046 279682 274102
rect 279738 274046 279808 274102
rect 279488 273978 279808 274046
rect 279488 273922 279558 273978
rect 279614 273922 279682 273978
rect 279738 273922 279808 273978
rect 279488 273888 279808 273922
rect 310208 274350 310528 274384
rect 310208 274294 310278 274350
rect 310334 274294 310402 274350
rect 310458 274294 310528 274350
rect 310208 274226 310528 274294
rect 310208 274170 310278 274226
rect 310334 274170 310402 274226
rect 310458 274170 310528 274226
rect 310208 274102 310528 274170
rect 310208 274046 310278 274102
rect 310334 274046 310402 274102
rect 310458 274046 310528 274102
rect 310208 273978 310528 274046
rect 310208 273922 310278 273978
rect 310334 273922 310402 273978
rect 310458 273922 310528 273978
rect 310208 273888 310528 273922
rect 340928 274350 341248 274384
rect 340928 274294 340998 274350
rect 341054 274294 341122 274350
rect 341178 274294 341248 274350
rect 340928 274226 341248 274294
rect 340928 274170 340998 274226
rect 341054 274170 341122 274226
rect 341178 274170 341248 274226
rect 340928 274102 341248 274170
rect 340928 274046 340998 274102
rect 341054 274046 341122 274102
rect 341178 274046 341248 274102
rect 340928 273978 341248 274046
rect 340928 273922 340998 273978
rect 341054 273922 341122 273978
rect 341178 273922 341248 273978
rect 340928 273888 341248 273922
rect 79808 262350 80128 262384
rect 79808 262294 79878 262350
rect 79934 262294 80002 262350
rect 80058 262294 80128 262350
rect 79808 262226 80128 262294
rect 79808 262170 79878 262226
rect 79934 262170 80002 262226
rect 80058 262170 80128 262226
rect 79808 262102 80128 262170
rect 79808 262046 79878 262102
rect 79934 262046 80002 262102
rect 80058 262046 80128 262102
rect 79808 261978 80128 262046
rect 79808 261922 79878 261978
rect 79934 261922 80002 261978
rect 80058 261922 80128 261978
rect 79808 261888 80128 261922
rect 110528 262350 110848 262384
rect 110528 262294 110598 262350
rect 110654 262294 110722 262350
rect 110778 262294 110848 262350
rect 110528 262226 110848 262294
rect 110528 262170 110598 262226
rect 110654 262170 110722 262226
rect 110778 262170 110848 262226
rect 110528 262102 110848 262170
rect 110528 262046 110598 262102
rect 110654 262046 110722 262102
rect 110778 262046 110848 262102
rect 110528 261978 110848 262046
rect 110528 261922 110598 261978
rect 110654 261922 110722 261978
rect 110778 261922 110848 261978
rect 110528 261888 110848 261922
rect 141248 262350 141568 262384
rect 141248 262294 141318 262350
rect 141374 262294 141442 262350
rect 141498 262294 141568 262350
rect 141248 262226 141568 262294
rect 141248 262170 141318 262226
rect 141374 262170 141442 262226
rect 141498 262170 141568 262226
rect 141248 262102 141568 262170
rect 141248 262046 141318 262102
rect 141374 262046 141442 262102
rect 141498 262046 141568 262102
rect 141248 261978 141568 262046
rect 141248 261922 141318 261978
rect 141374 261922 141442 261978
rect 141498 261922 141568 261978
rect 141248 261888 141568 261922
rect 171968 262350 172288 262384
rect 171968 262294 172038 262350
rect 172094 262294 172162 262350
rect 172218 262294 172288 262350
rect 171968 262226 172288 262294
rect 171968 262170 172038 262226
rect 172094 262170 172162 262226
rect 172218 262170 172288 262226
rect 171968 262102 172288 262170
rect 171968 262046 172038 262102
rect 172094 262046 172162 262102
rect 172218 262046 172288 262102
rect 171968 261978 172288 262046
rect 171968 261922 172038 261978
rect 172094 261922 172162 261978
rect 172218 261922 172288 261978
rect 171968 261888 172288 261922
rect 202688 262350 203008 262384
rect 202688 262294 202758 262350
rect 202814 262294 202882 262350
rect 202938 262294 203008 262350
rect 202688 262226 203008 262294
rect 202688 262170 202758 262226
rect 202814 262170 202882 262226
rect 202938 262170 203008 262226
rect 202688 262102 203008 262170
rect 202688 262046 202758 262102
rect 202814 262046 202882 262102
rect 202938 262046 203008 262102
rect 202688 261978 203008 262046
rect 202688 261922 202758 261978
rect 202814 261922 202882 261978
rect 202938 261922 203008 261978
rect 202688 261888 203008 261922
rect 233408 262350 233728 262384
rect 233408 262294 233478 262350
rect 233534 262294 233602 262350
rect 233658 262294 233728 262350
rect 233408 262226 233728 262294
rect 233408 262170 233478 262226
rect 233534 262170 233602 262226
rect 233658 262170 233728 262226
rect 233408 262102 233728 262170
rect 233408 262046 233478 262102
rect 233534 262046 233602 262102
rect 233658 262046 233728 262102
rect 233408 261978 233728 262046
rect 233408 261922 233478 261978
rect 233534 261922 233602 261978
rect 233658 261922 233728 261978
rect 233408 261888 233728 261922
rect 264128 262350 264448 262384
rect 264128 262294 264198 262350
rect 264254 262294 264322 262350
rect 264378 262294 264448 262350
rect 264128 262226 264448 262294
rect 264128 262170 264198 262226
rect 264254 262170 264322 262226
rect 264378 262170 264448 262226
rect 264128 262102 264448 262170
rect 264128 262046 264198 262102
rect 264254 262046 264322 262102
rect 264378 262046 264448 262102
rect 264128 261978 264448 262046
rect 264128 261922 264198 261978
rect 264254 261922 264322 261978
rect 264378 261922 264448 261978
rect 264128 261888 264448 261922
rect 294848 262350 295168 262384
rect 294848 262294 294918 262350
rect 294974 262294 295042 262350
rect 295098 262294 295168 262350
rect 294848 262226 295168 262294
rect 294848 262170 294918 262226
rect 294974 262170 295042 262226
rect 295098 262170 295168 262226
rect 294848 262102 295168 262170
rect 294848 262046 294918 262102
rect 294974 262046 295042 262102
rect 295098 262046 295168 262102
rect 294848 261978 295168 262046
rect 294848 261922 294918 261978
rect 294974 261922 295042 261978
rect 295098 261922 295168 261978
rect 294848 261888 295168 261922
rect 325568 262350 325888 262384
rect 325568 262294 325638 262350
rect 325694 262294 325762 262350
rect 325818 262294 325888 262350
rect 325568 262226 325888 262294
rect 325568 262170 325638 262226
rect 325694 262170 325762 262226
rect 325818 262170 325888 262226
rect 325568 262102 325888 262170
rect 325568 262046 325638 262102
rect 325694 262046 325762 262102
rect 325818 262046 325888 262102
rect 325568 261978 325888 262046
rect 325568 261922 325638 261978
rect 325694 261922 325762 261978
rect 325818 261922 325888 261978
rect 325568 261888 325888 261922
rect 348874 262350 349494 279922
rect 356288 280350 356608 280384
rect 356288 280294 356358 280350
rect 356414 280294 356482 280350
rect 356538 280294 356608 280350
rect 356288 280226 356608 280294
rect 356288 280170 356358 280226
rect 356414 280170 356482 280226
rect 356538 280170 356608 280226
rect 356288 280102 356608 280170
rect 356288 280046 356358 280102
rect 356414 280046 356482 280102
rect 356538 280046 356608 280102
rect 356288 279978 356608 280046
rect 356288 279922 356358 279978
rect 356414 279922 356482 279978
rect 356538 279922 356608 279978
rect 356288 279888 356608 279922
rect 363154 274350 363774 291922
rect 363154 274294 363250 274350
rect 363306 274294 363374 274350
rect 363430 274294 363498 274350
rect 363554 274294 363622 274350
rect 363678 274294 363774 274350
rect 363154 274226 363774 274294
rect 363154 274170 363250 274226
rect 363306 274170 363374 274226
rect 363430 274170 363498 274226
rect 363554 274170 363622 274226
rect 363678 274170 363774 274226
rect 363154 274102 363774 274170
rect 363154 274046 363250 274102
rect 363306 274046 363374 274102
rect 363430 274046 363498 274102
rect 363554 274046 363622 274102
rect 363678 274046 363774 274102
rect 363154 273978 363774 274046
rect 363154 273922 363250 273978
rect 363306 273922 363374 273978
rect 363430 273922 363498 273978
rect 363554 273922 363622 273978
rect 363678 273922 363774 273978
rect 348874 262294 348970 262350
rect 349026 262294 349094 262350
rect 349150 262294 349218 262350
rect 349274 262294 349342 262350
rect 349398 262294 349494 262350
rect 348874 262226 349494 262294
rect 348874 262170 348970 262226
rect 349026 262170 349094 262226
rect 349150 262170 349218 262226
rect 349274 262170 349342 262226
rect 349398 262170 349494 262226
rect 348874 262102 349494 262170
rect 348874 262046 348970 262102
rect 349026 262046 349094 262102
rect 349150 262046 349218 262102
rect 349274 262046 349342 262102
rect 349398 262046 349494 262102
rect 348874 261978 349494 262046
rect 348874 261922 348970 261978
rect 349026 261922 349094 261978
rect 349150 261922 349218 261978
rect 349274 261922 349342 261978
rect 349398 261922 349494 261978
rect 57154 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 57774 256350
rect 57154 256226 57774 256294
rect 57154 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 57774 256226
rect 57154 256102 57774 256170
rect 57154 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 57774 256102
rect 57154 255978 57774 256046
rect 57154 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 57774 255978
rect 57154 238350 57774 255922
rect 64448 256350 64768 256384
rect 64448 256294 64518 256350
rect 64574 256294 64642 256350
rect 64698 256294 64768 256350
rect 64448 256226 64768 256294
rect 64448 256170 64518 256226
rect 64574 256170 64642 256226
rect 64698 256170 64768 256226
rect 64448 256102 64768 256170
rect 64448 256046 64518 256102
rect 64574 256046 64642 256102
rect 64698 256046 64768 256102
rect 64448 255978 64768 256046
rect 64448 255922 64518 255978
rect 64574 255922 64642 255978
rect 64698 255922 64768 255978
rect 64448 255888 64768 255922
rect 95168 256350 95488 256384
rect 95168 256294 95238 256350
rect 95294 256294 95362 256350
rect 95418 256294 95488 256350
rect 95168 256226 95488 256294
rect 95168 256170 95238 256226
rect 95294 256170 95362 256226
rect 95418 256170 95488 256226
rect 95168 256102 95488 256170
rect 95168 256046 95238 256102
rect 95294 256046 95362 256102
rect 95418 256046 95488 256102
rect 95168 255978 95488 256046
rect 95168 255922 95238 255978
rect 95294 255922 95362 255978
rect 95418 255922 95488 255978
rect 95168 255888 95488 255922
rect 125888 256350 126208 256384
rect 125888 256294 125958 256350
rect 126014 256294 126082 256350
rect 126138 256294 126208 256350
rect 125888 256226 126208 256294
rect 125888 256170 125958 256226
rect 126014 256170 126082 256226
rect 126138 256170 126208 256226
rect 125888 256102 126208 256170
rect 125888 256046 125958 256102
rect 126014 256046 126082 256102
rect 126138 256046 126208 256102
rect 125888 255978 126208 256046
rect 125888 255922 125958 255978
rect 126014 255922 126082 255978
rect 126138 255922 126208 255978
rect 125888 255888 126208 255922
rect 156608 256350 156928 256384
rect 156608 256294 156678 256350
rect 156734 256294 156802 256350
rect 156858 256294 156928 256350
rect 156608 256226 156928 256294
rect 156608 256170 156678 256226
rect 156734 256170 156802 256226
rect 156858 256170 156928 256226
rect 156608 256102 156928 256170
rect 156608 256046 156678 256102
rect 156734 256046 156802 256102
rect 156858 256046 156928 256102
rect 156608 255978 156928 256046
rect 156608 255922 156678 255978
rect 156734 255922 156802 255978
rect 156858 255922 156928 255978
rect 156608 255888 156928 255922
rect 187328 256350 187648 256384
rect 187328 256294 187398 256350
rect 187454 256294 187522 256350
rect 187578 256294 187648 256350
rect 187328 256226 187648 256294
rect 187328 256170 187398 256226
rect 187454 256170 187522 256226
rect 187578 256170 187648 256226
rect 187328 256102 187648 256170
rect 187328 256046 187398 256102
rect 187454 256046 187522 256102
rect 187578 256046 187648 256102
rect 187328 255978 187648 256046
rect 187328 255922 187398 255978
rect 187454 255922 187522 255978
rect 187578 255922 187648 255978
rect 187328 255888 187648 255922
rect 218048 256350 218368 256384
rect 218048 256294 218118 256350
rect 218174 256294 218242 256350
rect 218298 256294 218368 256350
rect 218048 256226 218368 256294
rect 218048 256170 218118 256226
rect 218174 256170 218242 256226
rect 218298 256170 218368 256226
rect 218048 256102 218368 256170
rect 218048 256046 218118 256102
rect 218174 256046 218242 256102
rect 218298 256046 218368 256102
rect 218048 255978 218368 256046
rect 218048 255922 218118 255978
rect 218174 255922 218242 255978
rect 218298 255922 218368 255978
rect 218048 255888 218368 255922
rect 248768 256350 249088 256384
rect 248768 256294 248838 256350
rect 248894 256294 248962 256350
rect 249018 256294 249088 256350
rect 248768 256226 249088 256294
rect 248768 256170 248838 256226
rect 248894 256170 248962 256226
rect 249018 256170 249088 256226
rect 248768 256102 249088 256170
rect 248768 256046 248838 256102
rect 248894 256046 248962 256102
rect 249018 256046 249088 256102
rect 248768 255978 249088 256046
rect 248768 255922 248838 255978
rect 248894 255922 248962 255978
rect 249018 255922 249088 255978
rect 248768 255888 249088 255922
rect 279488 256350 279808 256384
rect 279488 256294 279558 256350
rect 279614 256294 279682 256350
rect 279738 256294 279808 256350
rect 279488 256226 279808 256294
rect 279488 256170 279558 256226
rect 279614 256170 279682 256226
rect 279738 256170 279808 256226
rect 279488 256102 279808 256170
rect 279488 256046 279558 256102
rect 279614 256046 279682 256102
rect 279738 256046 279808 256102
rect 279488 255978 279808 256046
rect 279488 255922 279558 255978
rect 279614 255922 279682 255978
rect 279738 255922 279808 255978
rect 279488 255888 279808 255922
rect 310208 256350 310528 256384
rect 310208 256294 310278 256350
rect 310334 256294 310402 256350
rect 310458 256294 310528 256350
rect 310208 256226 310528 256294
rect 310208 256170 310278 256226
rect 310334 256170 310402 256226
rect 310458 256170 310528 256226
rect 310208 256102 310528 256170
rect 310208 256046 310278 256102
rect 310334 256046 310402 256102
rect 310458 256046 310528 256102
rect 310208 255978 310528 256046
rect 310208 255922 310278 255978
rect 310334 255922 310402 255978
rect 310458 255922 310528 255978
rect 310208 255888 310528 255922
rect 340928 256350 341248 256384
rect 340928 256294 340998 256350
rect 341054 256294 341122 256350
rect 341178 256294 341248 256350
rect 340928 256226 341248 256294
rect 340928 256170 340998 256226
rect 341054 256170 341122 256226
rect 341178 256170 341248 256226
rect 340928 256102 341248 256170
rect 340928 256046 340998 256102
rect 341054 256046 341122 256102
rect 341178 256046 341248 256102
rect 340928 255978 341248 256046
rect 340928 255922 340998 255978
rect 341054 255922 341122 255978
rect 341178 255922 341248 255978
rect 340928 255888 341248 255922
rect 79808 244350 80128 244384
rect 79808 244294 79878 244350
rect 79934 244294 80002 244350
rect 80058 244294 80128 244350
rect 79808 244226 80128 244294
rect 79808 244170 79878 244226
rect 79934 244170 80002 244226
rect 80058 244170 80128 244226
rect 79808 244102 80128 244170
rect 79808 244046 79878 244102
rect 79934 244046 80002 244102
rect 80058 244046 80128 244102
rect 79808 243978 80128 244046
rect 79808 243922 79878 243978
rect 79934 243922 80002 243978
rect 80058 243922 80128 243978
rect 79808 243888 80128 243922
rect 110528 244350 110848 244384
rect 110528 244294 110598 244350
rect 110654 244294 110722 244350
rect 110778 244294 110848 244350
rect 110528 244226 110848 244294
rect 110528 244170 110598 244226
rect 110654 244170 110722 244226
rect 110778 244170 110848 244226
rect 110528 244102 110848 244170
rect 110528 244046 110598 244102
rect 110654 244046 110722 244102
rect 110778 244046 110848 244102
rect 110528 243978 110848 244046
rect 110528 243922 110598 243978
rect 110654 243922 110722 243978
rect 110778 243922 110848 243978
rect 110528 243888 110848 243922
rect 141248 244350 141568 244384
rect 141248 244294 141318 244350
rect 141374 244294 141442 244350
rect 141498 244294 141568 244350
rect 141248 244226 141568 244294
rect 141248 244170 141318 244226
rect 141374 244170 141442 244226
rect 141498 244170 141568 244226
rect 141248 244102 141568 244170
rect 141248 244046 141318 244102
rect 141374 244046 141442 244102
rect 141498 244046 141568 244102
rect 141248 243978 141568 244046
rect 141248 243922 141318 243978
rect 141374 243922 141442 243978
rect 141498 243922 141568 243978
rect 141248 243888 141568 243922
rect 171968 244350 172288 244384
rect 171968 244294 172038 244350
rect 172094 244294 172162 244350
rect 172218 244294 172288 244350
rect 171968 244226 172288 244294
rect 171968 244170 172038 244226
rect 172094 244170 172162 244226
rect 172218 244170 172288 244226
rect 171968 244102 172288 244170
rect 171968 244046 172038 244102
rect 172094 244046 172162 244102
rect 172218 244046 172288 244102
rect 171968 243978 172288 244046
rect 171968 243922 172038 243978
rect 172094 243922 172162 243978
rect 172218 243922 172288 243978
rect 171968 243888 172288 243922
rect 202688 244350 203008 244384
rect 202688 244294 202758 244350
rect 202814 244294 202882 244350
rect 202938 244294 203008 244350
rect 202688 244226 203008 244294
rect 202688 244170 202758 244226
rect 202814 244170 202882 244226
rect 202938 244170 203008 244226
rect 202688 244102 203008 244170
rect 202688 244046 202758 244102
rect 202814 244046 202882 244102
rect 202938 244046 203008 244102
rect 202688 243978 203008 244046
rect 202688 243922 202758 243978
rect 202814 243922 202882 243978
rect 202938 243922 203008 243978
rect 202688 243888 203008 243922
rect 233408 244350 233728 244384
rect 233408 244294 233478 244350
rect 233534 244294 233602 244350
rect 233658 244294 233728 244350
rect 233408 244226 233728 244294
rect 233408 244170 233478 244226
rect 233534 244170 233602 244226
rect 233658 244170 233728 244226
rect 233408 244102 233728 244170
rect 233408 244046 233478 244102
rect 233534 244046 233602 244102
rect 233658 244046 233728 244102
rect 233408 243978 233728 244046
rect 233408 243922 233478 243978
rect 233534 243922 233602 243978
rect 233658 243922 233728 243978
rect 233408 243888 233728 243922
rect 264128 244350 264448 244384
rect 264128 244294 264198 244350
rect 264254 244294 264322 244350
rect 264378 244294 264448 244350
rect 264128 244226 264448 244294
rect 264128 244170 264198 244226
rect 264254 244170 264322 244226
rect 264378 244170 264448 244226
rect 264128 244102 264448 244170
rect 264128 244046 264198 244102
rect 264254 244046 264322 244102
rect 264378 244046 264448 244102
rect 264128 243978 264448 244046
rect 264128 243922 264198 243978
rect 264254 243922 264322 243978
rect 264378 243922 264448 243978
rect 264128 243888 264448 243922
rect 294848 244350 295168 244384
rect 294848 244294 294918 244350
rect 294974 244294 295042 244350
rect 295098 244294 295168 244350
rect 294848 244226 295168 244294
rect 294848 244170 294918 244226
rect 294974 244170 295042 244226
rect 295098 244170 295168 244226
rect 294848 244102 295168 244170
rect 294848 244046 294918 244102
rect 294974 244046 295042 244102
rect 295098 244046 295168 244102
rect 294848 243978 295168 244046
rect 294848 243922 294918 243978
rect 294974 243922 295042 243978
rect 295098 243922 295168 243978
rect 294848 243888 295168 243922
rect 325568 244350 325888 244384
rect 325568 244294 325638 244350
rect 325694 244294 325762 244350
rect 325818 244294 325888 244350
rect 325568 244226 325888 244294
rect 325568 244170 325638 244226
rect 325694 244170 325762 244226
rect 325818 244170 325888 244226
rect 325568 244102 325888 244170
rect 325568 244046 325638 244102
rect 325694 244046 325762 244102
rect 325818 244046 325888 244102
rect 325568 243978 325888 244046
rect 325568 243922 325638 243978
rect 325694 243922 325762 243978
rect 325818 243922 325888 243978
rect 325568 243888 325888 243922
rect 348874 244350 349494 261922
rect 356288 262350 356608 262384
rect 356288 262294 356358 262350
rect 356414 262294 356482 262350
rect 356538 262294 356608 262350
rect 356288 262226 356608 262294
rect 356288 262170 356358 262226
rect 356414 262170 356482 262226
rect 356538 262170 356608 262226
rect 356288 262102 356608 262170
rect 356288 262046 356358 262102
rect 356414 262046 356482 262102
rect 356538 262046 356608 262102
rect 356288 261978 356608 262046
rect 356288 261922 356358 261978
rect 356414 261922 356482 261978
rect 356538 261922 356608 261978
rect 356288 261888 356608 261922
rect 363154 256350 363774 273922
rect 363154 256294 363250 256350
rect 363306 256294 363374 256350
rect 363430 256294 363498 256350
rect 363554 256294 363622 256350
rect 363678 256294 363774 256350
rect 363154 256226 363774 256294
rect 363154 256170 363250 256226
rect 363306 256170 363374 256226
rect 363430 256170 363498 256226
rect 363554 256170 363622 256226
rect 363678 256170 363774 256226
rect 363154 256102 363774 256170
rect 363154 256046 363250 256102
rect 363306 256046 363374 256102
rect 363430 256046 363498 256102
rect 363554 256046 363622 256102
rect 363678 256046 363774 256102
rect 363154 255978 363774 256046
rect 363154 255922 363250 255978
rect 363306 255922 363374 255978
rect 363430 255922 363498 255978
rect 363554 255922 363622 255978
rect 363678 255922 363774 255978
rect 348874 244294 348970 244350
rect 349026 244294 349094 244350
rect 349150 244294 349218 244350
rect 349274 244294 349342 244350
rect 349398 244294 349494 244350
rect 348874 244226 349494 244294
rect 348874 244170 348970 244226
rect 349026 244170 349094 244226
rect 349150 244170 349218 244226
rect 349274 244170 349342 244226
rect 349398 244170 349494 244226
rect 348874 244102 349494 244170
rect 348874 244046 348970 244102
rect 349026 244046 349094 244102
rect 349150 244046 349218 244102
rect 349274 244046 349342 244102
rect 349398 244046 349494 244102
rect 348874 243978 349494 244046
rect 348874 243922 348970 243978
rect 349026 243922 349094 243978
rect 349150 243922 349218 243978
rect 349274 243922 349342 243978
rect 349398 243922 349494 243978
rect 57154 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 57774 238350
rect 57154 238226 57774 238294
rect 57154 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 57774 238226
rect 57154 238102 57774 238170
rect 57154 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 57774 238102
rect 57154 237978 57774 238046
rect 57154 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 57774 237978
rect 57154 220350 57774 237922
rect 64448 238350 64768 238384
rect 64448 238294 64518 238350
rect 64574 238294 64642 238350
rect 64698 238294 64768 238350
rect 64448 238226 64768 238294
rect 64448 238170 64518 238226
rect 64574 238170 64642 238226
rect 64698 238170 64768 238226
rect 64448 238102 64768 238170
rect 64448 238046 64518 238102
rect 64574 238046 64642 238102
rect 64698 238046 64768 238102
rect 64448 237978 64768 238046
rect 64448 237922 64518 237978
rect 64574 237922 64642 237978
rect 64698 237922 64768 237978
rect 64448 237888 64768 237922
rect 95168 238350 95488 238384
rect 95168 238294 95238 238350
rect 95294 238294 95362 238350
rect 95418 238294 95488 238350
rect 95168 238226 95488 238294
rect 95168 238170 95238 238226
rect 95294 238170 95362 238226
rect 95418 238170 95488 238226
rect 95168 238102 95488 238170
rect 95168 238046 95238 238102
rect 95294 238046 95362 238102
rect 95418 238046 95488 238102
rect 95168 237978 95488 238046
rect 95168 237922 95238 237978
rect 95294 237922 95362 237978
rect 95418 237922 95488 237978
rect 95168 237888 95488 237922
rect 125888 238350 126208 238384
rect 125888 238294 125958 238350
rect 126014 238294 126082 238350
rect 126138 238294 126208 238350
rect 125888 238226 126208 238294
rect 125888 238170 125958 238226
rect 126014 238170 126082 238226
rect 126138 238170 126208 238226
rect 125888 238102 126208 238170
rect 125888 238046 125958 238102
rect 126014 238046 126082 238102
rect 126138 238046 126208 238102
rect 125888 237978 126208 238046
rect 125888 237922 125958 237978
rect 126014 237922 126082 237978
rect 126138 237922 126208 237978
rect 125888 237888 126208 237922
rect 156608 238350 156928 238384
rect 156608 238294 156678 238350
rect 156734 238294 156802 238350
rect 156858 238294 156928 238350
rect 156608 238226 156928 238294
rect 156608 238170 156678 238226
rect 156734 238170 156802 238226
rect 156858 238170 156928 238226
rect 156608 238102 156928 238170
rect 156608 238046 156678 238102
rect 156734 238046 156802 238102
rect 156858 238046 156928 238102
rect 156608 237978 156928 238046
rect 156608 237922 156678 237978
rect 156734 237922 156802 237978
rect 156858 237922 156928 237978
rect 156608 237888 156928 237922
rect 187328 238350 187648 238384
rect 187328 238294 187398 238350
rect 187454 238294 187522 238350
rect 187578 238294 187648 238350
rect 187328 238226 187648 238294
rect 187328 238170 187398 238226
rect 187454 238170 187522 238226
rect 187578 238170 187648 238226
rect 187328 238102 187648 238170
rect 187328 238046 187398 238102
rect 187454 238046 187522 238102
rect 187578 238046 187648 238102
rect 187328 237978 187648 238046
rect 187328 237922 187398 237978
rect 187454 237922 187522 237978
rect 187578 237922 187648 237978
rect 187328 237888 187648 237922
rect 218048 238350 218368 238384
rect 218048 238294 218118 238350
rect 218174 238294 218242 238350
rect 218298 238294 218368 238350
rect 218048 238226 218368 238294
rect 218048 238170 218118 238226
rect 218174 238170 218242 238226
rect 218298 238170 218368 238226
rect 218048 238102 218368 238170
rect 218048 238046 218118 238102
rect 218174 238046 218242 238102
rect 218298 238046 218368 238102
rect 218048 237978 218368 238046
rect 218048 237922 218118 237978
rect 218174 237922 218242 237978
rect 218298 237922 218368 237978
rect 218048 237888 218368 237922
rect 248768 238350 249088 238384
rect 248768 238294 248838 238350
rect 248894 238294 248962 238350
rect 249018 238294 249088 238350
rect 248768 238226 249088 238294
rect 248768 238170 248838 238226
rect 248894 238170 248962 238226
rect 249018 238170 249088 238226
rect 248768 238102 249088 238170
rect 248768 238046 248838 238102
rect 248894 238046 248962 238102
rect 249018 238046 249088 238102
rect 248768 237978 249088 238046
rect 248768 237922 248838 237978
rect 248894 237922 248962 237978
rect 249018 237922 249088 237978
rect 248768 237888 249088 237922
rect 279488 238350 279808 238384
rect 279488 238294 279558 238350
rect 279614 238294 279682 238350
rect 279738 238294 279808 238350
rect 279488 238226 279808 238294
rect 279488 238170 279558 238226
rect 279614 238170 279682 238226
rect 279738 238170 279808 238226
rect 279488 238102 279808 238170
rect 279488 238046 279558 238102
rect 279614 238046 279682 238102
rect 279738 238046 279808 238102
rect 279488 237978 279808 238046
rect 279488 237922 279558 237978
rect 279614 237922 279682 237978
rect 279738 237922 279808 237978
rect 279488 237888 279808 237922
rect 310208 238350 310528 238384
rect 310208 238294 310278 238350
rect 310334 238294 310402 238350
rect 310458 238294 310528 238350
rect 310208 238226 310528 238294
rect 310208 238170 310278 238226
rect 310334 238170 310402 238226
rect 310458 238170 310528 238226
rect 310208 238102 310528 238170
rect 310208 238046 310278 238102
rect 310334 238046 310402 238102
rect 310458 238046 310528 238102
rect 310208 237978 310528 238046
rect 310208 237922 310278 237978
rect 310334 237922 310402 237978
rect 310458 237922 310528 237978
rect 310208 237888 310528 237922
rect 340928 238350 341248 238384
rect 340928 238294 340998 238350
rect 341054 238294 341122 238350
rect 341178 238294 341248 238350
rect 340928 238226 341248 238294
rect 340928 238170 340998 238226
rect 341054 238170 341122 238226
rect 341178 238170 341248 238226
rect 340928 238102 341248 238170
rect 340928 238046 340998 238102
rect 341054 238046 341122 238102
rect 341178 238046 341248 238102
rect 340928 237978 341248 238046
rect 340928 237922 340998 237978
rect 341054 237922 341122 237978
rect 341178 237922 341248 237978
rect 340928 237888 341248 237922
rect 79808 226350 80128 226384
rect 79808 226294 79878 226350
rect 79934 226294 80002 226350
rect 80058 226294 80128 226350
rect 79808 226226 80128 226294
rect 79808 226170 79878 226226
rect 79934 226170 80002 226226
rect 80058 226170 80128 226226
rect 79808 226102 80128 226170
rect 79808 226046 79878 226102
rect 79934 226046 80002 226102
rect 80058 226046 80128 226102
rect 79808 225978 80128 226046
rect 79808 225922 79878 225978
rect 79934 225922 80002 225978
rect 80058 225922 80128 225978
rect 79808 225888 80128 225922
rect 110528 226350 110848 226384
rect 110528 226294 110598 226350
rect 110654 226294 110722 226350
rect 110778 226294 110848 226350
rect 110528 226226 110848 226294
rect 110528 226170 110598 226226
rect 110654 226170 110722 226226
rect 110778 226170 110848 226226
rect 110528 226102 110848 226170
rect 110528 226046 110598 226102
rect 110654 226046 110722 226102
rect 110778 226046 110848 226102
rect 110528 225978 110848 226046
rect 110528 225922 110598 225978
rect 110654 225922 110722 225978
rect 110778 225922 110848 225978
rect 110528 225888 110848 225922
rect 141248 226350 141568 226384
rect 141248 226294 141318 226350
rect 141374 226294 141442 226350
rect 141498 226294 141568 226350
rect 141248 226226 141568 226294
rect 141248 226170 141318 226226
rect 141374 226170 141442 226226
rect 141498 226170 141568 226226
rect 141248 226102 141568 226170
rect 141248 226046 141318 226102
rect 141374 226046 141442 226102
rect 141498 226046 141568 226102
rect 141248 225978 141568 226046
rect 141248 225922 141318 225978
rect 141374 225922 141442 225978
rect 141498 225922 141568 225978
rect 141248 225888 141568 225922
rect 171968 226350 172288 226384
rect 171968 226294 172038 226350
rect 172094 226294 172162 226350
rect 172218 226294 172288 226350
rect 171968 226226 172288 226294
rect 171968 226170 172038 226226
rect 172094 226170 172162 226226
rect 172218 226170 172288 226226
rect 171968 226102 172288 226170
rect 171968 226046 172038 226102
rect 172094 226046 172162 226102
rect 172218 226046 172288 226102
rect 171968 225978 172288 226046
rect 171968 225922 172038 225978
rect 172094 225922 172162 225978
rect 172218 225922 172288 225978
rect 171968 225888 172288 225922
rect 202688 226350 203008 226384
rect 202688 226294 202758 226350
rect 202814 226294 202882 226350
rect 202938 226294 203008 226350
rect 202688 226226 203008 226294
rect 202688 226170 202758 226226
rect 202814 226170 202882 226226
rect 202938 226170 203008 226226
rect 202688 226102 203008 226170
rect 202688 226046 202758 226102
rect 202814 226046 202882 226102
rect 202938 226046 203008 226102
rect 202688 225978 203008 226046
rect 202688 225922 202758 225978
rect 202814 225922 202882 225978
rect 202938 225922 203008 225978
rect 202688 225888 203008 225922
rect 233408 226350 233728 226384
rect 233408 226294 233478 226350
rect 233534 226294 233602 226350
rect 233658 226294 233728 226350
rect 233408 226226 233728 226294
rect 233408 226170 233478 226226
rect 233534 226170 233602 226226
rect 233658 226170 233728 226226
rect 233408 226102 233728 226170
rect 233408 226046 233478 226102
rect 233534 226046 233602 226102
rect 233658 226046 233728 226102
rect 233408 225978 233728 226046
rect 233408 225922 233478 225978
rect 233534 225922 233602 225978
rect 233658 225922 233728 225978
rect 233408 225888 233728 225922
rect 264128 226350 264448 226384
rect 264128 226294 264198 226350
rect 264254 226294 264322 226350
rect 264378 226294 264448 226350
rect 264128 226226 264448 226294
rect 264128 226170 264198 226226
rect 264254 226170 264322 226226
rect 264378 226170 264448 226226
rect 264128 226102 264448 226170
rect 264128 226046 264198 226102
rect 264254 226046 264322 226102
rect 264378 226046 264448 226102
rect 264128 225978 264448 226046
rect 264128 225922 264198 225978
rect 264254 225922 264322 225978
rect 264378 225922 264448 225978
rect 264128 225888 264448 225922
rect 294848 226350 295168 226384
rect 294848 226294 294918 226350
rect 294974 226294 295042 226350
rect 295098 226294 295168 226350
rect 294848 226226 295168 226294
rect 294848 226170 294918 226226
rect 294974 226170 295042 226226
rect 295098 226170 295168 226226
rect 294848 226102 295168 226170
rect 294848 226046 294918 226102
rect 294974 226046 295042 226102
rect 295098 226046 295168 226102
rect 294848 225978 295168 226046
rect 294848 225922 294918 225978
rect 294974 225922 295042 225978
rect 295098 225922 295168 225978
rect 294848 225888 295168 225922
rect 325568 226350 325888 226384
rect 325568 226294 325638 226350
rect 325694 226294 325762 226350
rect 325818 226294 325888 226350
rect 325568 226226 325888 226294
rect 325568 226170 325638 226226
rect 325694 226170 325762 226226
rect 325818 226170 325888 226226
rect 325568 226102 325888 226170
rect 325568 226046 325638 226102
rect 325694 226046 325762 226102
rect 325818 226046 325888 226102
rect 325568 225978 325888 226046
rect 325568 225922 325638 225978
rect 325694 225922 325762 225978
rect 325818 225922 325888 225978
rect 325568 225888 325888 225922
rect 348874 226350 349494 243922
rect 356288 244350 356608 244384
rect 356288 244294 356358 244350
rect 356414 244294 356482 244350
rect 356538 244294 356608 244350
rect 356288 244226 356608 244294
rect 356288 244170 356358 244226
rect 356414 244170 356482 244226
rect 356538 244170 356608 244226
rect 356288 244102 356608 244170
rect 356288 244046 356358 244102
rect 356414 244046 356482 244102
rect 356538 244046 356608 244102
rect 356288 243978 356608 244046
rect 356288 243922 356358 243978
rect 356414 243922 356482 243978
rect 356538 243922 356608 243978
rect 356288 243888 356608 243922
rect 363154 238350 363774 255922
rect 363154 238294 363250 238350
rect 363306 238294 363374 238350
rect 363430 238294 363498 238350
rect 363554 238294 363622 238350
rect 363678 238294 363774 238350
rect 363154 238226 363774 238294
rect 363154 238170 363250 238226
rect 363306 238170 363374 238226
rect 363430 238170 363498 238226
rect 363554 238170 363622 238226
rect 363678 238170 363774 238226
rect 363154 238102 363774 238170
rect 363154 238046 363250 238102
rect 363306 238046 363374 238102
rect 363430 238046 363498 238102
rect 363554 238046 363622 238102
rect 363678 238046 363774 238102
rect 363154 237978 363774 238046
rect 363154 237922 363250 237978
rect 363306 237922 363374 237978
rect 363430 237922 363498 237978
rect 363554 237922 363622 237978
rect 363678 237922 363774 237978
rect 348874 226294 348970 226350
rect 349026 226294 349094 226350
rect 349150 226294 349218 226350
rect 349274 226294 349342 226350
rect 349398 226294 349494 226350
rect 348874 226226 349494 226294
rect 348874 226170 348970 226226
rect 349026 226170 349094 226226
rect 349150 226170 349218 226226
rect 349274 226170 349342 226226
rect 349398 226170 349494 226226
rect 348874 226102 349494 226170
rect 348874 226046 348970 226102
rect 349026 226046 349094 226102
rect 349150 226046 349218 226102
rect 349274 226046 349342 226102
rect 349398 226046 349494 226102
rect 348874 225978 349494 226046
rect 348874 225922 348970 225978
rect 349026 225922 349094 225978
rect 349150 225922 349218 225978
rect 349274 225922 349342 225978
rect 349398 225922 349494 225978
rect 57154 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 57774 220350
rect 57154 220226 57774 220294
rect 57154 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 57774 220226
rect 57154 220102 57774 220170
rect 57154 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 57774 220102
rect 57154 219978 57774 220046
rect 57154 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 57774 219978
rect 57154 202350 57774 219922
rect 64448 220350 64768 220384
rect 64448 220294 64518 220350
rect 64574 220294 64642 220350
rect 64698 220294 64768 220350
rect 64448 220226 64768 220294
rect 64448 220170 64518 220226
rect 64574 220170 64642 220226
rect 64698 220170 64768 220226
rect 64448 220102 64768 220170
rect 64448 220046 64518 220102
rect 64574 220046 64642 220102
rect 64698 220046 64768 220102
rect 64448 219978 64768 220046
rect 64448 219922 64518 219978
rect 64574 219922 64642 219978
rect 64698 219922 64768 219978
rect 64448 219888 64768 219922
rect 95168 220350 95488 220384
rect 95168 220294 95238 220350
rect 95294 220294 95362 220350
rect 95418 220294 95488 220350
rect 95168 220226 95488 220294
rect 95168 220170 95238 220226
rect 95294 220170 95362 220226
rect 95418 220170 95488 220226
rect 95168 220102 95488 220170
rect 95168 220046 95238 220102
rect 95294 220046 95362 220102
rect 95418 220046 95488 220102
rect 95168 219978 95488 220046
rect 95168 219922 95238 219978
rect 95294 219922 95362 219978
rect 95418 219922 95488 219978
rect 95168 219888 95488 219922
rect 125888 220350 126208 220384
rect 125888 220294 125958 220350
rect 126014 220294 126082 220350
rect 126138 220294 126208 220350
rect 125888 220226 126208 220294
rect 125888 220170 125958 220226
rect 126014 220170 126082 220226
rect 126138 220170 126208 220226
rect 125888 220102 126208 220170
rect 125888 220046 125958 220102
rect 126014 220046 126082 220102
rect 126138 220046 126208 220102
rect 125888 219978 126208 220046
rect 125888 219922 125958 219978
rect 126014 219922 126082 219978
rect 126138 219922 126208 219978
rect 125888 219888 126208 219922
rect 156608 220350 156928 220384
rect 156608 220294 156678 220350
rect 156734 220294 156802 220350
rect 156858 220294 156928 220350
rect 156608 220226 156928 220294
rect 156608 220170 156678 220226
rect 156734 220170 156802 220226
rect 156858 220170 156928 220226
rect 156608 220102 156928 220170
rect 156608 220046 156678 220102
rect 156734 220046 156802 220102
rect 156858 220046 156928 220102
rect 156608 219978 156928 220046
rect 156608 219922 156678 219978
rect 156734 219922 156802 219978
rect 156858 219922 156928 219978
rect 156608 219888 156928 219922
rect 187328 220350 187648 220384
rect 187328 220294 187398 220350
rect 187454 220294 187522 220350
rect 187578 220294 187648 220350
rect 187328 220226 187648 220294
rect 187328 220170 187398 220226
rect 187454 220170 187522 220226
rect 187578 220170 187648 220226
rect 187328 220102 187648 220170
rect 187328 220046 187398 220102
rect 187454 220046 187522 220102
rect 187578 220046 187648 220102
rect 187328 219978 187648 220046
rect 187328 219922 187398 219978
rect 187454 219922 187522 219978
rect 187578 219922 187648 219978
rect 187328 219888 187648 219922
rect 218048 220350 218368 220384
rect 218048 220294 218118 220350
rect 218174 220294 218242 220350
rect 218298 220294 218368 220350
rect 218048 220226 218368 220294
rect 218048 220170 218118 220226
rect 218174 220170 218242 220226
rect 218298 220170 218368 220226
rect 218048 220102 218368 220170
rect 218048 220046 218118 220102
rect 218174 220046 218242 220102
rect 218298 220046 218368 220102
rect 218048 219978 218368 220046
rect 218048 219922 218118 219978
rect 218174 219922 218242 219978
rect 218298 219922 218368 219978
rect 218048 219888 218368 219922
rect 248768 220350 249088 220384
rect 248768 220294 248838 220350
rect 248894 220294 248962 220350
rect 249018 220294 249088 220350
rect 248768 220226 249088 220294
rect 248768 220170 248838 220226
rect 248894 220170 248962 220226
rect 249018 220170 249088 220226
rect 248768 220102 249088 220170
rect 248768 220046 248838 220102
rect 248894 220046 248962 220102
rect 249018 220046 249088 220102
rect 248768 219978 249088 220046
rect 248768 219922 248838 219978
rect 248894 219922 248962 219978
rect 249018 219922 249088 219978
rect 248768 219888 249088 219922
rect 279488 220350 279808 220384
rect 279488 220294 279558 220350
rect 279614 220294 279682 220350
rect 279738 220294 279808 220350
rect 279488 220226 279808 220294
rect 279488 220170 279558 220226
rect 279614 220170 279682 220226
rect 279738 220170 279808 220226
rect 279488 220102 279808 220170
rect 279488 220046 279558 220102
rect 279614 220046 279682 220102
rect 279738 220046 279808 220102
rect 279488 219978 279808 220046
rect 279488 219922 279558 219978
rect 279614 219922 279682 219978
rect 279738 219922 279808 219978
rect 279488 219888 279808 219922
rect 310208 220350 310528 220384
rect 310208 220294 310278 220350
rect 310334 220294 310402 220350
rect 310458 220294 310528 220350
rect 310208 220226 310528 220294
rect 310208 220170 310278 220226
rect 310334 220170 310402 220226
rect 310458 220170 310528 220226
rect 310208 220102 310528 220170
rect 310208 220046 310278 220102
rect 310334 220046 310402 220102
rect 310458 220046 310528 220102
rect 310208 219978 310528 220046
rect 310208 219922 310278 219978
rect 310334 219922 310402 219978
rect 310458 219922 310528 219978
rect 310208 219888 310528 219922
rect 340928 220350 341248 220384
rect 340928 220294 340998 220350
rect 341054 220294 341122 220350
rect 341178 220294 341248 220350
rect 340928 220226 341248 220294
rect 340928 220170 340998 220226
rect 341054 220170 341122 220226
rect 341178 220170 341248 220226
rect 340928 220102 341248 220170
rect 340928 220046 340998 220102
rect 341054 220046 341122 220102
rect 341178 220046 341248 220102
rect 340928 219978 341248 220046
rect 340928 219922 340998 219978
rect 341054 219922 341122 219978
rect 341178 219922 341248 219978
rect 340928 219888 341248 219922
rect 79808 208350 80128 208384
rect 79808 208294 79878 208350
rect 79934 208294 80002 208350
rect 80058 208294 80128 208350
rect 79808 208226 80128 208294
rect 79808 208170 79878 208226
rect 79934 208170 80002 208226
rect 80058 208170 80128 208226
rect 79808 208102 80128 208170
rect 79808 208046 79878 208102
rect 79934 208046 80002 208102
rect 80058 208046 80128 208102
rect 79808 207978 80128 208046
rect 79808 207922 79878 207978
rect 79934 207922 80002 207978
rect 80058 207922 80128 207978
rect 79808 207888 80128 207922
rect 110528 208350 110848 208384
rect 110528 208294 110598 208350
rect 110654 208294 110722 208350
rect 110778 208294 110848 208350
rect 110528 208226 110848 208294
rect 110528 208170 110598 208226
rect 110654 208170 110722 208226
rect 110778 208170 110848 208226
rect 110528 208102 110848 208170
rect 110528 208046 110598 208102
rect 110654 208046 110722 208102
rect 110778 208046 110848 208102
rect 110528 207978 110848 208046
rect 110528 207922 110598 207978
rect 110654 207922 110722 207978
rect 110778 207922 110848 207978
rect 110528 207888 110848 207922
rect 141248 208350 141568 208384
rect 141248 208294 141318 208350
rect 141374 208294 141442 208350
rect 141498 208294 141568 208350
rect 141248 208226 141568 208294
rect 141248 208170 141318 208226
rect 141374 208170 141442 208226
rect 141498 208170 141568 208226
rect 141248 208102 141568 208170
rect 141248 208046 141318 208102
rect 141374 208046 141442 208102
rect 141498 208046 141568 208102
rect 141248 207978 141568 208046
rect 141248 207922 141318 207978
rect 141374 207922 141442 207978
rect 141498 207922 141568 207978
rect 141248 207888 141568 207922
rect 171968 208350 172288 208384
rect 171968 208294 172038 208350
rect 172094 208294 172162 208350
rect 172218 208294 172288 208350
rect 171968 208226 172288 208294
rect 171968 208170 172038 208226
rect 172094 208170 172162 208226
rect 172218 208170 172288 208226
rect 171968 208102 172288 208170
rect 171968 208046 172038 208102
rect 172094 208046 172162 208102
rect 172218 208046 172288 208102
rect 171968 207978 172288 208046
rect 171968 207922 172038 207978
rect 172094 207922 172162 207978
rect 172218 207922 172288 207978
rect 171968 207888 172288 207922
rect 202688 208350 203008 208384
rect 202688 208294 202758 208350
rect 202814 208294 202882 208350
rect 202938 208294 203008 208350
rect 202688 208226 203008 208294
rect 202688 208170 202758 208226
rect 202814 208170 202882 208226
rect 202938 208170 203008 208226
rect 202688 208102 203008 208170
rect 202688 208046 202758 208102
rect 202814 208046 202882 208102
rect 202938 208046 203008 208102
rect 202688 207978 203008 208046
rect 202688 207922 202758 207978
rect 202814 207922 202882 207978
rect 202938 207922 203008 207978
rect 202688 207888 203008 207922
rect 233408 208350 233728 208384
rect 233408 208294 233478 208350
rect 233534 208294 233602 208350
rect 233658 208294 233728 208350
rect 233408 208226 233728 208294
rect 233408 208170 233478 208226
rect 233534 208170 233602 208226
rect 233658 208170 233728 208226
rect 233408 208102 233728 208170
rect 233408 208046 233478 208102
rect 233534 208046 233602 208102
rect 233658 208046 233728 208102
rect 233408 207978 233728 208046
rect 233408 207922 233478 207978
rect 233534 207922 233602 207978
rect 233658 207922 233728 207978
rect 233408 207888 233728 207922
rect 264128 208350 264448 208384
rect 264128 208294 264198 208350
rect 264254 208294 264322 208350
rect 264378 208294 264448 208350
rect 264128 208226 264448 208294
rect 264128 208170 264198 208226
rect 264254 208170 264322 208226
rect 264378 208170 264448 208226
rect 264128 208102 264448 208170
rect 264128 208046 264198 208102
rect 264254 208046 264322 208102
rect 264378 208046 264448 208102
rect 264128 207978 264448 208046
rect 264128 207922 264198 207978
rect 264254 207922 264322 207978
rect 264378 207922 264448 207978
rect 264128 207888 264448 207922
rect 294848 208350 295168 208384
rect 294848 208294 294918 208350
rect 294974 208294 295042 208350
rect 295098 208294 295168 208350
rect 294848 208226 295168 208294
rect 294848 208170 294918 208226
rect 294974 208170 295042 208226
rect 295098 208170 295168 208226
rect 294848 208102 295168 208170
rect 294848 208046 294918 208102
rect 294974 208046 295042 208102
rect 295098 208046 295168 208102
rect 294848 207978 295168 208046
rect 294848 207922 294918 207978
rect 294974 207922 295042 207978
rect 295098 207922 295168 207978
rect 294848 207888 295168 207922
rect 325568 208350 325888 208384
rect 325568 208294 325638 208350
rect 325694 208294 325762 208350
rect 325818 208294 325888 208350
rect 325568 208226 325888 208294
rect 325568 208170 325638 208226
rect 325694 208170 325762 208226
rect 325818 208170 325888 208226
rect 325568 208102 325888 208170
rect 325568 208046 325638 208102
rect 325694 208046 325762 208102
rect 325818 208046 325888 208102
rect 325568 207978 325888 208046
rect 325568 207922 325638 207978
rect 325694 207922 325762 207978
rect 325818 207922 325888 207978
rect 325568 207888 325888 207922
rect 348874 208350 349494 225922
rect 356288 226350 356608 226384
rect 356288 226294 356358 226350
rect 356414 226294 356482 226350
rect 356538 226294 356608 226350
rect 356288 226226 356608 226294
rect 356288 226170 356358 226226
rect 356414 226170 356482 226226
rect 356538 226170 356608 226226
rect 356288 226102 356608 226170
rect 356288 226046 356358 226102
rect 356414 226046 356482 226102
rect 356538 226046 356608 226102
rect 356288 225978 356608 226046
rect 356288 225922 356358 225978
rect 356414 225922 356482 225978
rect 356538 225922 356608 225978
rect 356288 225888 356608 225922
rect 363154 220350 363774 237922
rect 363154 220294 363250 220350
rect 363306 220294 363374 220350
rect 363430 220294 363498 220350
rect 363554 220294 363622 220350
rect 363678 220294 363774 220350
rect 363154 220226 363774 220294
rect 363154 220170 363250 220226
rect 363306 220170 363374 220226
rect 363430 220170 363498 220226
rect 363554 220170 363622 220226
rect 363678 220170 363774 220226
rect 363154 220102 363774 220170
rect 363154 220046 363250 220102
rect 363306 220046 363374 220102
rect 363430 220046 363498 220102
rect 363554 220046 363622 220102
rect 363678 220046 363774 220102
rect 363154 219978 363774 220046
rect 363154 219922 363250 219978
rect 363306 219922 363374 219978
rect 363430 219922 363498 219978
rect 363554 219922 363622 219978
rect 363678 219922 363774 219978
rect 348874 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 349494 208350
rect 348874 208226 349494 208294
rect 348874 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 349494 208226
rect 348874 208102 349494 208170
rect 348874 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 349494 208102
rect 348874 207978 349494 208046
rect 348874 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 349494 207978
rect 57154 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 57774 202350
rect 57154 202226 57774 202294
rect 57154 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 57774 202226
rect 57154 202102 57774 202170
rect 57154 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 57774 202102
rect 57154 201978 57774 202046
rect 57154 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 57774 201978
rect 57154 184350 57774 201922
rect 64448 202350 64768 202384
rect 64448 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 64768 202350
rect 64448 202226 64768 202294
rect 64448 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 64768 202226
rect 64448 202102 64768 202170
rect 64448 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 64768 202102
rect 64448 201978 64768 202046
rect 64448 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 64768 201978
rect 64448 201888 64768 201922
rect 95168 202350 95488 202384
rect 95168 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 95488 202350
rect 95168 202226 95488 202294
rect 95168 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 95488 202226
rect 95168 202102 95488 202170
rect 95168 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 95488 202102
rect 95168 201978 95488 202046
rect 95168 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 95488 201978
rect 95168 201888 95488 201922
rect 125888 202350 126208 202384
rect 125888 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 126208 202350
rect 125888 202226 126208 202294
rect 125888 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 126208 202226
rect 125888 202102 126208 202170
rect 125888 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 126208 202102
rect 125888 201978 126208 202046
rect 125888 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 126208 201978
rect 125888 201888 126208 201922
rect 156608 202350 156928 202384
rect 156608 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 156928 202350
rect 156608 202226 156928 202294
rect 156608 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 156928 202226
rect 156608 202102 156928 202170
rect 156608 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 156928 202102
rect 156608 201978 156928 202046
rect 156608 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 156928 201978
rect 156608 201888 156928 201922
rect 187328 202350 187648 202384
rect 187328 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 187648 202350
rect 187328 202226 187648 202294
rect 187328 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 187648 202226
rect 187328 202102 187648 202170
rect 187328 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 187648 202102
rect 187328 201978 187648 202046
rect 187328 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 187648 201978
rect 187328 201888 187648 201922
rect 218048 202350 218368 202384
rect 218048 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 218368 202350
rect 218048 202226 218368 202294
rect 218048 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 218368 202226
rect 218048 202102 218368 202170
rect 218048 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 218368 202102
rect 218048 201978 218368 202046
rect 218048 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 218368 201978
rect 218048 201888 218368 201922
rect 248768 202350 249088 202384
rect 248768 202294 248838 202350
rect 248894 202294 248962 202350
rect 249018 202294 249088 202350
rect 248768 202226 249088 202294
rect 248768 202170 248838 202226
rect 248894 202170 248962 202226
rect 249018 202170 249088 202226
rect 248768 202102 249088 202170
rect 248768 202046 248838 202102
rect 248894 202046 248962 202102
rect 249018 202046 249088 202102
rect 248768 201978 249088 202046
rect 248768 201922 248838 201978
rect 248894 201922 248962 201978
rect 249018 201922 249088 201978
rect 248768 201888 249088 201922
rect 279488 202350 279808 202384
rect 279488 202294 279558 202350
rect 279614 202294 279682 202350
rect 279738 202294 279808 202350
rect 279488 202226 279808 202294
rect 279488 202170 279558 202226
rect 279614 202170 279682 202226
rect 279738 202170 279808 202226
rect 279488 202102 279808 202170
rect 279488 202046 279558 202102
rect 279614 202046 279682 202102
rect 279738 202046 279808 202102
rect 279488 201978 279808 202046
rect 279488 201922 279558 201978
rect 279614 201922 279682 201978
rect 279738 201922 279808 201978
rect 279488 201888 279808 201922
rect 310208 202350 310528 202384
rect 310208 202294 310278 202350
rect 310334 202294 310402 202350
rect 310458 202294 310528 202350
rect 310208 202226 310528 202294
rect 310208 202170 310278 202226
rect 310334 202170 310402 202226
rect 310458 202170 310528 202226
rect 310208 202102 310528 202170
rect 310208 202046 310278 202102
rect 310334 202046 310402 202102
rect 310458 202046 310528 202102
rect 310208 201978 310528 202046
rect 310208 201922 310278 201978
rect 310334 201922 310402 201978
rect 310458 201922 310528 201978
rect 310208 201888 310528 201922
rect 340928 202350 341248 202384
rect 340928 202294 340998 202350
rect 341054 202294 341122 202350
rect 341178 202294 341248 202350
rect 340928 202226 341248 202294
rect 340928 202170 340998 202226
rect 341054 202170 341122 202226
rect 341178 202170 341248 202226
rect 340928 202102 341248 202170
rect 340928 202046 340998 202102
rect 341054 202046 341122 202102
rect 341178 202046 341248 202102
rect 340928 201978 341248 202046
rect 340928 201922 340998 201978
rect 341054 201922 341122 201978
rect 341178 201922 341248 201978
rect 340928 201888 341248 201922
rect 79808 190350 80128 190384
rect 79808 190294 79878 190350
rect 79934 190294 80002 190350
rect 80058 190294 80128 190350
rect 79808 190226 80128 190294
rect 79808 190170 79878 190226
rect 79934 190170 80002 190226
rect 80058 190170 80128 190226
rect 79808 190102 80128 190170
rect 79808 190046 79878 190102
rect 79934 190046 80002 190102
rect 80058 190046 80128 190102
rect 79808 189978 80128 190046
rect 79808 189922 79878 189978
rect 79934 189922 80002 189978
rect 80058 189922 80128 189978
rect 79808 189888 80128 189922
rect 110528 190350 110848 190384
rect 110528 190294 110598 190350
rect 110654 190294 110722 190350
rect 110778 190294 110848 190350
rect 110528 190226 110848 190294
rect 110528 190170 110598 190226
rect 110654 190170 110722 190226
rect 110778 190170 110848 190226
rect 110528 190102 110848 190170
rect 110528 190046 110598 190102
rect 110654 190046 110722 190102
rect 110778 190046 110848 190102
rect 110528 189978 110848 190046
rect 110528 189922 110598 189978
rect 110654 189922 110722 189978
rect 110778 189922 110848 189978
rect 110528 189888 110848 189922
rect 141248 190350 141568 190384
rect 141248 190294 141318 190350
rect 141374 190294 141442 190350
rect 141498 190294 141568 190350
rect 141248 190226 141568 190294
rect 141248 190170 141318 190226
rect 141374 190170 141442 190226
rect 141498 190170 141568 190226
rect 141248 190102 141568 190170
rect 141248 190046 141318 190102
rect 141374 190046 141442 190102
rect 141498 190046 141568 190102
rect 141248 189978 141568 190046
rect 141248 189922 141318 189978
rect 141374 189922 141442 189978
rect 141498 189922 141568 189978
rect 141248 189888 141568 189922
rect 171968 190350 172288 190384
rect 171968 190294 172038 190350
rect 172094 190294 172162 190350
rect 172218 190294 172288 190350
rect 171968 190226 172288 190294
rect 171968 190170 172038 190226
rect 172094 190170 172162 190226
rect 172218 190170 172288 190226
rect 171968 190102 172288 190170
rect 171968 190046 172038 190102
rect 172094 190046 172162 190102
rect 172218 190046 172288 190102
rect 171968 189978 172288 190046
rect 171968 189922 172038 189978
rect 172094 189922 172162 189978
rect 172218 189922 172288 189978
rect 171968 189888 172288 189922
rect 202688 190350 203008 190384
rect 202688 190294 202758 190350
rect 202814 190294 202882 190350
rect 202938 190294 203008 190350
rect 202688 190226 203008 190294
rect 202688 190170 202758 190226
rect 202814 190170 202882 190226
rect 202938 190170 203008 190226
rect 202688 190102 203008 190170
rect 202688 190046 202758 190102
rect 202814 190046 202882 190102
rect 202938 190046 203008 190102
rect 202688 189978 203008 190046
rect 202688 189922 202758 189978
rect 202814 189922 202882 189978
rect 202938 189922 203008 189978
rect 202688 189888 203008 189922
rect 233408 190350 233728 190384
rect 233408 190294 233478 190350
rect 233534 190294 233602 190350
rect 233658 190294 233728 190350
rect 233408 190226 233728 190294
rect 233408 190170 233478 190226
rect 233534 190170 233602 190226
rect 233658 190170 233728 190226
rect 233408 190102 233728 190170
rect 233408 190046 233478 190102
rect 233534 190046 233602 190102
rect 233658 190046 233728 190102
rect 233408 189978 233728 190046
rect 233408 189922 233478 189978
rect 233534 189922 233602 189978
rect 233658 189922 233728 189978
rect 233408 189888 233728 189922
rect 264128 190350 264448 190384
rect 264128 190294 264198 190350
rect 264254 190294 264322 190350
rect 264378 190294 264448 190350
rect 264128 190226 264448 190294
rect 264128 190170 264198 190226
rect 264254 190170 264322 190226
rect 264378 190170 264448 190226
rect 264128 190102 264448 190170
rect 264128 190046 264198 190102
rect 264254 190046 264322 190102
rect 264378 190046 264448 190102
rect 264128 189978 264448 190046
rect 264128 189922 264198 189978
rect 264254 189922 264322 189978
rect 264378 189922 264448 189978
rect 264128 189888 264448 189922
rect 294848 190350 295168 190384
rect 294848 190294 294918 190350
rect 294974 190294 295042 190350
rect 295098 190294 295168 190350
rect 294848 190226 295168 190294
rect 294848 190170 294918 190226
rect 294974 190170 295042 190226
rect 295098 190170 295168 190226
rect 294848 190102 295168 190170
rect 294848 190046 294918 190102
rect 294974 190046 295042 190102
rect 295098 190046 295168 190102
rect 294848 189978 295168 190046
rect 294848 189922 294918 189978
rect 294974 189922 295042 189978
rect 295098 189922 295168 189978
rect 294848 189888 295168 189922
rect 325568 190350 325888 190384
rect 325568 190294 325638 190350
rect 325694 190294 325762 190350
rect 325818 190294 325888 190350
rect 325568 190226 325888 190294
rect 325568 190170 325638 190226
rect 325694 190170 325762 190226
rect 325818 190170 325888 190226
rect 325568 190102 325888 190170
rect 325568 190046 325638 190102
rect 325694 190046 325762 190102
rect 325818 190046 325888 190102
rect 325568 189978 325888 190046
rect 325568 189922 325638 189978
rect 325694 189922 325762 189978
rect 325818 189922 325888 189978
rect 325568 189888 325888 189922
rect 348874 190350 349494 207922
rect 356288 208350 356608 208384
rect 356288 208294 356358 208350
rect 356414 208294 356482 208350
rect 356538 208294 356608 208350
rect 356288 208226 356608 208294
rect 356288 208170 356358 208226
rect 356414 208170 356482 208226
rect 356538 208170 356608 208226
rect 356288 208102 356608 208170
rect 356288 208046 356358 208102
rect 356414 208046 356482 208102
rect 356538 208046 356608 208102
rect 356288 207978 356608 208046
rect 356288 207922 356358 207978
rect 356414 207922 356482 207978
rect 356538 207922 356608 207978
rect 356288 207888 356608 207922
rect 363154 202350 363774 219922
rect 363154 202294 363250 202350
rect 363306 202294 363374 202350
rect 363430 202294 363498 202350
rect 363554 202294 363622 202350
rect 363678 202294 363774 202350
rect 363154 202226 363774 202294
rect 363154 202170 363250 202226
rect 363306 202170 363374 202226
rect 363430 202170 363498 202226
rect 363554 202170 363622 202226
rect 363678 202170 363774 202226
rect 363154 202102 363774 202170
rect 363154 202046 363250 202102
rect 363306 202046 363374 202102
rect 363430 202046 363498 202102
rect 363554 202046 363622 202102
rect 363678 202046 363774 202102
rect 363154 201978 363774 202046
rect 363154 201922 363250 201978
rect 363306 201922 363374 201978
rect 363430 201922 363498 201978
rect 363554 201922 363622 201978
rect 363678 201922 363774 201978
rect 348874 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 349494 190350
rect 348874 190226 349494 190294
rect 348874 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 349494 190226
rect 348874 190102 349494 190170
rect 348874 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 349494 190102
rect 348874 189978 349494 190046
rect 348874 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 349494 189978
rect 57154 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 57774 184350
rect 57154 184226 57774 184294
rect 57154 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 57774 184226
rect 57154 184102 57774 184170
rect 57154 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 57774 184102
rect 57154 183978 57774 184046
rect 57154 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 57774 183978
rect 57154 166350 57774 183922
rect 64448 184350 64768 184384
rect 64448 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 64768 184350
rect 64448 184226 64768 184294
rect 64448 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 64768 184226
rect 64448 184102 64768 184170
rect 64448 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 64768 184102
rect 64448 183978 64768 184046
rect 64448 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 64768 183978
rect 64448 183888 64768 183922
rect 95168 184350 95488 184384
rect 95168 184294 95238 184350
rect 95294 184294 95362 184350
rect 95418 184294 95488 184350
rect 95168 184226 95488 184294
rect 95168 184170 95238 184226
rect 95294 184170 95362 184226
rect 95418 184170 95488 184226
rect 95168 184102 95488 184170
rect 95168 184046 95238 184102
rect 95294 184046 95362 184102
rect 95418 184046 95488 184102
rect 95168 183978 95488 184046
rect 95168 183922 95238 183978
rect 95294 183922 95362 183978
rect 95418 183922 95488 183978
rect 95168 183888 95488 183922
rect 125888 184350 126208 184384
rect 125888 184294 125958 184350
rect 126014 184294 126082 184350
rect 126138 184294 126208 184350
rect 125888 184226 126208 184294
rect 125888 184170 125958 184226
rect 126014 184170 126082 184226
rect 126138 184170 126208 184226
rect 125888 184102 126208 184170
rect 125888 184046 125958 184102
rect 126014 184046 126082 184102
rect 126138 184046 126208 184102
rect 125888 183978 126208 184046
rect 125888 183922 125958 183978
rect 126014 183922 126082 183978
rect 126138 183922 126208 183978
rect 125888 183888 126208 183922
rect 156608 184350 156928 184384
rect 156608 184294 156678 184350
rect 156734 184294 156802 184350
rect 156858 184294 156928 184350
rect 156608 184226 156928 184294
rect 156608 184170 156678 184226
rect 156734 184170 156802 184226
rect 156858 184170 156928 184226
rect 156608 184102 156928 184170
rect 156608 184046 156678 184102
rect 156734 184046 156802 184102
rect 156858 184046 156928 184102
rect 156608 183978 156928 184046
rect 156608 183922 156678 183978
rect 156734 183922 156802 183978
rect 156858 183922 156928 183978
rect 156608 183888 156928 183922
rect 187328 184350 187648 184384
rect 187328 184294 187398 184350
rect 187454 184294 187522 184350
rect 187578 184294 187648 184350
rect 187328 184226 187648 184294
rect 187328 184170 187398 184226
rect 187454 184170 187522 184226
rect 187578 184170 187648 184226
rect 187328 184102 187648 184170
rect 187328 184046 187398 184102
rect 187454 184046 187522 184102
rect 187578 184046 187648 184102
rect 187328 183978 187648 184046
rect 187328 183922 187398 183978
rect 187454 183922 187522 183978
rect 187578 183922 187648 183978
rect 187328 183888 187648 183922
rect 218048 184350 218368 184384
rect 218048 184294 218118 184350
rect 218174 184294 218242 184350
rect 218298 184294 218368 184350
rect 218048 184226 218368 184294
rect 218048 184170 218118 184226
rect 218174 184170 218242 184226
rect 218298 184170 218368 184226
rect 218048 184102 218368 184170
rect 218048 184046 218118 184102
rect 218174 184046 218242 184102
rect 218298 184046 218368 184102
rect 218048 183978 218368 184046
rect 218048 183922 218118 183978
rect 218174 183922 218242 183978
rect 218298 183922 218368 183978
rect 218048 183888 218368 183922
rect 248768 184350 249088 184384
rect 248768 184294 248838 184350
rect 248894 184294 248962 184350
rect 249018 184294 249088 184350
rect 248768 184226 249088 184294
rect 248768 184170 248838 184226
rect 248894 184170 248962 184226
rect 249018 184170 249088 184226
rect 248768 184102 249088 184170
rect 248768 184046 248838 184102
rect 248894 184046 248962 184102
rect 249018 184046 249088 184102
rect 248768 183978 249088 184046
rect 248768 183922 248838 183978
rect 248894 183922 248962 183978
rect 249018 183922 249088 183978
rect 248768 183888 249088 183922
rect 279488 184350 279808 184384
rect 279488 184294 279558 184350
rect 279614 184294 279682 184350
rect 279738 184294 279808 184350
rect 279488 184226 279808 184294
rect 279488 184170 279558 184226
rect 279614 184170 279682 184226
rect 279738 184170 279808 184226
rect 279488 184102 279808 184170
rect 279488 184046 279558 184102
rect 279614 184046 279682 184102
rect 279738 184046 279808 184102
rect 279488 183978 279808 184046
rect 279488 183922 279558 183978
rect 279614 183922 279682 183978
rect 279738 183922 279808 183978
rect 279488 183888 279808 183922
rect 310208 184350 310528 184384
rect 310208 184294 310278 184350
rect 310334 184294 310402 184350
rect 310458 184294 310528 184350
rect 310208 184226 310528 184294
rect 310208 184170 310278 184226
rect 310334 184170 310402 184226
rect 310458 184170 310528 184226
rect 310208 184102 310528 184170
rect 310208 184046 310278 184102
rect 310334 184046 310402 184102
rect 310458 184046 310528 184102
rect 310208 183978 310528 184046
rect 310208 183922 310278 183978
rect 310334 183922 310402 183978
rect 310458 183922 310528 183978
rect 310208 183888 310528 183922
rect 340928 184350 341248 184384
rect 340928 184294 340998 184350
rect 341054 184294 341122 184350
rect 341178 184294 341248 184350
rect 340928 184226 341248 184294
rect 340928 184170 340998 184226
rect 341054 184170 341122 184226
rect 341178 184170 341248 184226
rect 340928 184102 341248 184170
rect 340928 184046 340998 184102
rect 341054 184046 341122 184102
rect 341178 184046 341248 184102
rect 340928 183978 341248 184046
rect 340928 183922 340998 183978
rect 341054 183922 341122 183978
rect 341178 183922 341248 183978
rect 340928 183888 341248 183922
rect 79808 172350 80128 172384
rect 79808 172294 79878 172350
rect 79934 172294 80002 172350
rect 80058 172294 80128 172350
rect 79808 172226 80128 172294
rect 79808 172170 79878 172226
rect 79934 172170 80002 172226
rect 80058 172170 80128 172226
rect 79808 172102 80128 172170
rect 79808 172046 79878 172102
rect 79934 172046 80002 172102
rect 80058 172046 80128 172102
rect 79808 171978 80128 172046
rect 79808 171922 79878 171978
rect 79934 171922 80002 171978
rect 80058 171922 80128 171978
rect 79808 171888 80128 171922
rect 110528 172350 110848 172384
rect 110528 172294 110598 172350
rect 110654 172294 110722 172350
rect 110778 172294 110848 172350
rect 110528 172226 110848 172294
rect 110528 172170 110598 172226
rect 110654 172170 110722 172226
rect 110778 172170 110848 172226
rect 110528 172102 110848 172170
rect 110528 172046 110598 172102
rect 110654 172046 110722 172102
rect 110778 172046 110848 172102
rect 110528 171978 110848 172046
rect 110528 171922 110598 171978
rect 110654 171922 110722 171978
rect 110778 171922 110848 171978
rect 110528 171888 110848 171922
rect 141248 172350 141568 172384
rect 141248 172294 141318 172350
rect 141374 172294 141442 172350
rect 141498 172294 141568 172350
rect 141248 172226 141568 172294
rect 141248 172170 141318 172226
rect 141374 172170 141442 172226
rect 141498 172170 141568 172226
rect 141248 172102 141568 172170
rect 141248 172046 141318 172102
rect 141374 172046 141442 172102
rect 141498 172046 141568 172102
rect 141248 171978 141568 172046
rect 141248 171922 141318 171978
rect 141374 171922 141442 171978
rect 141498 171922 141568 171978
rect 141248 171888 141568 171922
rect 171968 172350 172288 172384
rect 171968 172294 172038 172350
rect 172094 172294 172162 172350
rect 172218 172294 172288 172350
rect 171968 172226 172288 172294
rect 171968 172170 172038 172226
rect 172094 172170 172162 172226
rect 172218 172170 172288 172226
rect 171968 172102 172288 172170
rect 171968 172046 172038 172102
rect 172094 172046 172162 172102
rect 172218 172046 172288 172102
rect 171968 171978 172288 172046
rect 171968 171922 172038 171978
rect 172094 171922 172162 171978
rect 172218 171922 172288 171978
rect 171968 171888 172288 171922
rect 202688 172350 203008 172384
rect 202688 172294 202758 172350
rect 202814 172294 202882 172350
rect 202938 172294 203008 172350
rect 202688 172226 203008 172294
rect 202688 172170 202758 172226
rect 202814 172170 202882 172226
rect 202938 172170 203008 172226
rect 202688 172102 203008 172170
rect 202688 172046 202758 172102
rect 202814 172046 202882 172102
rect 202938 172046 203008 172102
rect 202688 171978 203008 172046
rect 202688 171922 202758 171978
rect 202814 171922 202882 171978
rect 202938 171922 203008 171978
rect 202688 171888 203008 171922
rect 233408 172350 233728 172384
rect 233408 172294 233478 172350
rect 233534 172294 233602 172350
rect 233658 172294 233728 172350
rect 233408 172226 233728 172294
rect 233408 172170 233478 172226
rect 233534 172170 233602 172226
rect 233658 172170 233728 172226
rect 233408 172102 233728 172170
rect 233408 172046 233478 172102
rect 233534 172046 233602 172102
rect 233658 172046 233728 172102
rect 233408 171978 233728 172046
rect 233408 171922 233478 171978
rect 233534 171922 233602 171978
rect 233658 171922 233728 171978
rect 233408 171888 233728 171922
rect 264128 172350 264448 172384
rect 264128 172294 264198 172350
rect 264254 172294 264322 172350
rect 264378 172294 264448 172350
rect 264128 172226 264448 172294
rect 264128 172170 264198 172226
rect 264254 172170 264322 172226
rect 264378 172170 264448 172226
rect 264128 172102 264448 172170
rect 264128 172046 264198 172102
rect 264254 172046 264322 172102
rect 264378 172046 264448 172102
rect 264128 171978 264448 172046
rect 264128 171922 264198 171978
rect 264254 171922 264322 171978
rect 264378 171922 264448 171978
rect 264128 171888 264448 171922
rect 294848 172350 295168 172384
rect 294848 172294 294918 172350
rect 294974 172294 295042 172350
rect 295098 172294 295168 172350
rect 294848 172226 295168 172294
rect 294848 172170 294918 172226
rect 294974 172170 295042 172226
rect 295098 172170 295168 172226
rect 294848 172102 295168 172170
rect 294848 172046 294918 172102
rect 294974 172046 295042 172102
rect 295098 172046 295168 172102
rect 294848 171978 295168 172046
rect 294848 171922 294918 171978
rect 294974 171922 295042 171978
rect 295098 171922 295168 171978
rect 294848 171888 295168 171922
rect 325568 172350 325888 172384
rect 325568 172294 325638 172350
rect 325694 172294 325762 172350
rect 325818 172294 325888 172350
rect 325568 172226 325888 172294
rect 325568 172170 325638 172226
rect 325694 172170 325762 172226
rect 325818 172170 325888 172226
rect 325568 172102 325888 172170
rect 325568 172046 325638 172102
rect 325694 172046 325762 172102
rect 325818 172046 325888 172102
rect 325568 171978 325888 172046
rect 325568 171922 325638 171978
rect 325694 171922 325762 171978
rect 325818 171922 325888 171978
rect 325568 171888 325888 171922
rect 348874 172350 349494 189922
rect 356288 190350 356608 190384
rect 356288 190294 356358 190350
rect 356414 190294 356482 190350
rect 356538 190294 356608 190350
rect 356288 190226 356608 190294
rect 356288 190170 356358 190226
rect 356414 190170 356482 190226
rect 356538 190170 356608 190226
rect 356288 190102 356608 190170
rect 356288 190046 356358 190102
rect 356414 190046 356482 190102
rect 356538 190046 356608 190102
rect 356288 189978 356608 190046
rect 356288 189922 356358 189978
rect 356414 189922 356482 189978
rect 356538 189922 356608 189978
rect 356288 189888 356608 189922
rect 363154 184350 363774 201922
rect 363154 184294 363250 184350
rect 363306 184294 363374 184350
rect 363430 184294 363498 184350
rect 363554 184294 363622 184350
rect 363678 184294 363774 184350
rect 363154 184226 363774 184294
rect 363154 184170 363250 184226
rect 363306 184170 363374 184226
rect 363430 184170 363498 184226
rect 363554 184170 363622 184226
rect 363678 184170 363774 184226
rect 363154 184102 363774 184170
rect 363154 184046 363250 184102
rect 363306 184046 363374 184102
rect 363430 184046 363498 184102
rect 363554 184046 363622 184102
rect 363678 184046 363774 184102
rect 363154 183978 363774 184046
rect 363154 183922 363250 183978
rect 363306 183922 363374 183978
rect 363430 183922 363498 183978
rect 363554 183922 363622 183978
rect 363678 183922 363774 183978
rect 348874 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 349494 172350
rect 348874 172226 349494 172294
rect 348874 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 349494 172226
rect 348874 172102 349494 172170
rect 348874 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 349494 172102
rect 348874 171978 349494 172046
rect 348874 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 349494 171978
rect 57154 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 57774 166350
rect 57154 166226 57774 166294
rect 57154 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 57774 166226
rect 57154 166102 57774 166170
rect 57154 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 57774 166102
rect 57154 165978 57774 166046
rect 57154 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 57774 165978
rect 57154 148350 57774 165922
rect 64448 166350 64768 166384
rect 64448 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 64768 166350
rect 64448 166226 64768 166294
rect 64448 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 64768 166226
rect 64448 166102 64768 166170
rect 64448 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 64768 166102
rect 64448 165978 64768 166046
rect 64448 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 64768 165978
rect 64448 165888 64768 165922
rect 95168 166350 95488 166384
rect 95168 166294 95238 166350
rect 95294 166294 95362 166350
rect 95418 166294 95488 166350
rect 95168 166226 95488 166294
rect 95168 166170 95238 166226
rect 95294 166170 95362 166226
rect 95418 166170 95488 166226
rect 95168 166102 95488 166170
rect 95168 166046 95238 166102
rect 95294 166046 95362 166102
rect 95418 166046 95488 166102
rect 95168 165978 95488 166046
rect 95168 165922 95238 165978
rect 95294 165922 95362 165978
rect 95418 165922 95488 165978
rect 95168 165888 95488 165922
rect 125888 166350 126208 166384
rect 125888 166294 125958 166350
rect 126014 166294 126082 166350
rect 126138 166294 126208 166350
rect 125888 166226 126208 166294
rect 125888 166170 125958 166226
rect 126014 166170 126082 166226
rect 126138 166170 126208 166226
rect 125888 166102 126208 166170
rect 125888 166046 125958 166102
rect 126014 166046 126082 166102
rect 126138 166046 126208 166102
rect 125888 165978 126208 166046
rect 125888 165922 125958 165978
rect 126014 165922 126082 165978
rect 126138 165922 126208 165978
rect 125888 165888 126208 165922
rect 156608 166350 156928 166384
rect 156608 166294 156678 166350
rect 156734 166294 156802 166350
rect 156858 166294 156928 166350
rect 156608 166226 156928 166294
rect 156608 166170 156678 166226
rect 156734 166170 156802 166226
rect 156858 166170 156928 166226
rect 156608 166102 156928 166170
rect 156608 166046 156678 166102
rect 156734 166046 156802 166102
rect 156858 166046 156928 166102
rect 156608 165978 156928 166046
rect 156608 165922 156678 165978
rect 156734 165922 156802 165978
rect 156858 165922 156928 165978
rect 156608 165888 156928 165922
rect 187328 166350 187648 166384
rect 187328 166294 187398 166350
rect 187454 166294 187522 166350
rect 187578 166294 187648 166350
rect 187328 166226 187648 166294
rect 187328 166170 187398 166226
rect 187454 166170 187522 166226
rect 187578 166170 187648 166226
rect 187328 166102 187648 166170
rect 187328 166046 187398 166102
rect 187454 166046 187522 166102
rect 187578 166046 187648 166102
rect 187328 165978 187648 166046
rect 187328 165922 187398 165978
rect 187454 165922 187522 165978
rect 187578 165922 187648 165978
rect 187328 165888 187648 165922
rect 218048 166350 218368 166384
rect 218048 166294 218118 166350
rect 218174 166294 218242 166350
rect 218298 166294 218368 166350
rect 218048 166226 218368 166294
rect 218048 166170 218118 166226
rect 218174 166170 218242 166226
rect 218298 166170 218368 166226
rect 218048 166102 218368 166170
rect 218048 166046 218118 166102
rect 218174 166046 218242 166102
rect 218298 166046 218368 166102
rect 218048 165978 218368 166046
rect 218048 165922 218118 165978
rect 218174 165922 218242 165978
rect 218298 165922 218368 165978
rect 218048 165888 218368 165922
rect 248768 166350 249088 166384
rect 248768 166294 248838 166350
rect 248894 166294 248962 166350
rect 249018 166294 249088 166350
rect 248768 166226 249088 166294
rect 248768 166170 248838 166226
rect 248894 166170 248962 166226
rect 249018 166170 249088 166226
rect 248768 166102 249088 166170
rect 248768 166046 248838 166102
rect 248894 166046 248962 166102
rect 249018 166046 249088 166102
rect 248768 165978 249088 166046
rect 248768 165922 248838 165978
rect 248894 165922 248962 165978
rect 249018 165922 249088 165978
rect 248768 165888 249088 165922
rect 279488 166350 279808 166384
rect 279488 166294 279558 166350
rect 279614 166294 279682 166350
rect 279738 166294 279808 166350
rect 279488 166226 279808 166294
rect 279488 166170 279558 166226
rect 279614 166170 279682 166226
rect 279738 166170 279808 166226
rect 279488 166102 279808 166170
rect 279488 166046 279558 166102
rect 279614 166046 279682 166102
rect 279738 166046 279808 166102
rect 279488 165978 279808 166046
rect 279488 165922 279558 165978
rect 279614 165922 279682 165978
rect 279738 165922 279808 165978
rect 279488 165888 279808 165922
rect 310208 166350 310528 166384
rect 310208 166294 310278 166350
rect 310334 166294 310402 166350
rect 310458 166294 310528 166350
rect 310208 166226 310528 166294
rect 310208 166170 310278 166226
rect 310334 166170 310402 166226
rect 310458 166170 310528 166226
rect 310208 166102 310528 166170
rect 310208 166046 310278 166102
rect 310334 166046 310402 166102
rect 310458 166046 310528 166102
rect 310208 165978 310528 166046
rect 310208 165922 310278 165978
rect 310334 165922 310402 165978
rect 310458 165922 310528 165978
rect 310208 165888 310528 165922
rect 340928 166350 341248 166384
rect 340928 166294 340998 166350
rect 341054 166294 341122 166350
rect 341178 166294 341248 166350
rect 340928 166226 341248 166294
rect 340928 166170 340998 166226
rect 341054 166170 341122 166226
rect 341178 166170 341248 166226
rect 340928 166102 341248 166170
rect 340928 166046 340998 166102
rect 341054 166046 341122 166102
rect 341178 166046 341248 166102
rect 340928 165978 341248 166046
rect 340928 165922 340998 165978
rect 341054 165922 341122 165978
rect 341178 165922 341248 165978
rect 340928 165888 341248 165922
rect 79808 154350 80128 154384
rect 79808 154294 79878 154350
rect 79934 154294 80002 154350
rect 80058 154294 80128 154350
rect 79808 154226 80128 154294
rect 79808 154170 79878 154226
rect 79934 154170 80002 154226
rect 80058 154170 80128 154226
rect 79808 154102 80128 154170
rect 79808 154046 79878 154102
rect 79934 154046 80002 154102
rect 80058 154046 80128 154102
rect 79808 153978 80128 154046
rect 79808 153922 79878 153978
rect 79934 153922 80002 153978
rect 80058 153922 80128 153978
rect 79808 153888 80128 153922
rect 110528 154350 110848 154384
rect 110528 154294 110598 154350
rect 110654 154294 110722 154350
rect 110778 154294 110848 154350
rect 110528 154226 110848 154294
rect 110528 154170 110598 154226
rect 110654 154170 110722 154226
rect 110778 154170 110848 154226
rect 110528 154102 110848 154170
rect 110528 154046 110598 154102
rect 110654 154046 110722 154102
rect 110778 154046 110848 154102
rect 110528 153978 110848 154046
rect 110528 153922 110598 153978
rect 110654 153922 110722 153978
rect 110778 153922 110848 153978
rect 110528 153888 110848 153922
rect 141248 154350 141568 154384
rect 141248 154294 141318 154350
rect 141374 154294 141442 154350
rect 141498 154294 141568 154350
rect 141248 154226 141568 154294
rect 141248 154170 141318 154226
rect 141374 154170 141442 154226
rect 141498 154170 141568 154226
rect 141248 154102 141568 154170
rect 141248 154046 141318 154102
rect 141374 154046 141442 154102
rect 141498 154046 141568 154102
rect 141248 153978 141568 154046
rect 141248 153922 141318 153978
rect 141374 153922 141442 153978
rect 141498 153922 141568 153978
rect 141248 153888 141568 153922
rect 171968 154350 172288 154384
rect 171968 154294 172038 154350
rect 172094 154294 172162 154350
rect 172218 154294 172288 154350
rect 171968 154226 172288 154294
rect 171968 154170 172038 154226
rect 172094 154170 172162 154226
rect 172218 154170 172288 154226
rect 171968 154102 172288 154170
rect 171968 154046 172038 154102
rect 172094 154046 172162 154102
rect 172218 154046 172288 154102
rect 171968 153978 172288 154046
rect 171968 153922 172038 153978
rect 172094 153922 172162 153978
rect 172218 153922 172288 153978
rect 171968 153888 172288 153922
rect 202688 154350 203008 154384
rect 202688 154294 202758 154350
rect 202814 154294 202882 154350
rect 202938 154294 203008 154350
rect 202688 154226 203008 154294
rect 202688 154170 202758 154226
rect 202814 154170 202882 154226
rect 202938 154170 203008 154226
rect 202688 154102 203008 154170
rect 202688 154046 202758 154102
rect 202814 154046 202882 154102
rect 202938 154046 203008 154102
rect 202688 153978 203008 154046
rect 202688 153922 202758 153978
rect 202814 153922 202882 153978
rect 202938 153922 203008 153978
rect 202688 153888 203008 153922
rect 233408 154350 233728 154384
rect 233408 154294 233478 154350
rect 233534 154294 233602 154350
rect 233658 154294 233728 154350
rect 233408 154226 233728 154294
rect 233408 154170 233478 154226
rect 233534 154170 233602 154226
rect 233658 154170 233728 154226
rect 233408 154102 233728 154170
rect 233408 154046 233478 154102
rect 233534 154046 233602 154102
rect 233658 154046 233728 154102
rect 233408 153978 233728 154046
rect 233408 153922 233478 153978
rect 233534 153922 233602 153978
rect 233658 153922 233728 153978
rect 233408 153888 233728 153922
rect 264128 154350 264448 154384
rect 264128 154294 264198 154350
rect 264254 154294 264322 154350
rect 264378 154294 264448 154350
rect 264128 154226 264448 154294
rect 264128 154170 264198 154226
rect 264254 154170 264322 154226
rect 264378 154170 264448 154226
rect 264128 154102 264448 154170
rect 264128 154046 264198 154102
rect 264254 154046 264322 154102
rect 264378 154046 264448 154102
rect 264128 153978 264448 154046
rect 264128 153922 264198 153978
rect 264254 153922 264322 153978
rect 264378 153922 264448 153978
rect 264128 153888 264448 153922
rect 294848 154350 295168 154384
rect 294848 154294 294918 154350
rect 294974 154294 295042 154350
rect 295098 154294 295168 154350
rect 294848 154226 295168 154294
rect 294848 154170 294918 154226
rect 294974 154170 295042 154226
rect 295098 154170 295168 154226
rect 294848 154102 295168 154170
rect 294848 154046 294918 154102
rect 294974 154046 295042 154102
rect 295098 154046 295168 154102
rect 294848 153978 295168 154046
rect 294848 153922 294918 153978
rect 294974 153922 295042 153978
rect 295098 153922 295168 153978
rect 294848 153888 295168 153922
rect 325568 154350 325888 154384
rect 325568 154294 325638 154350
rect 325694 154294 325762 154350
rect 325818 154294 325888 154350
rect 325568 154226 325888 154294
rect 325568 154170 325638 154226
rect 325694 154170 325762 154226
rect 325818 154170 325888 154226
rect 325568 154102 325888 154170
rect 325568 154046 325638 154102
rect 325694 154046 325762 154102
rect 325818 154046 325888 154102
rect 325568 153978 325888 154046
rect 325568 153922 325638 153978
rect 325694 153922 325762 153978
rect 325818 153922 325888 153978
rect 325568 153888 325888 153922
rect 348874 154350 349494 171922
rect 356288 172350 356608 172384
rect 356288 172294 356358 172350
rect 356414 172294 356482 172350
rect 356538 172294 356608 172350
rect 356288 172226 356608 172294
rect 356288 172170 356358 172226
rect 356414 172170 356482 172226
rect 356538 172170 356608 172226
rect 356288 172102 356608 172170
rect 356288 172046 356358 172102
rect 356414 172046 356482 172102
rect 356538 172046 356608 172102
rect 356288 171978 356608 172046
rect 356288 171922 356358 171978
rect 356414 171922 356482 171978
rect 356538 171922 356608 171978
rect 356288 171888 356608 171922
rect 363154 166350 363774 183922
rect 363154 166294 363250 166350
rect 363306 166294 363374 166350
rect 363430 166294 363498 166350
rect 363554 166294 363622 166350
rect 363678 166294 363774 166350
rect 363154 166226 363774 166294
rect 363154 166170 363250 166226
rect 363306 166170 363374 166226
rect 363430 166170 363498 166226
rect 363554 166170 363622 166226
rect 363678 166170 363774 166226
rect 363154 166102 363774 166170
rect 363154 166046 363250 166102
rect 363306 166046 363374 166102
rect 363430 166046 363498 166102
rect 363554 166046 363622 166102
rect 363678 166046 363774 166102
rect 363154 165978 363774 166046
rect 363154 165922 363250 165978
rect 363306 165922 363374 165978
rect 363430 165922 363498 165978
rect 363554 165922 363622 165978
rect 363678 165922 363774 165978
rect 348874 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 349494 154350
rect 348874 154226 349494 154294
rect 348874 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 349494 154226
rect 348874 154102 349494 154170
rect 348874 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 349494 154102
rect 348874 153978 349494 154046
rect 348874 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 349494 153978
rect 57154 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 57774 148350
rect 57154 148226 57774 148294
rect 57154 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 57774 148226
rect 57154 148102 57774 148170
rect 57154 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 57774 148102
rect 57154 147978 57774 148046
rect 57154 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 57774 147978
rect 57154 130350 57774 147922
rect 64448 148350 64768 148384
rect 64448 148294 64518 148350
rect 64574 148294 64642 148350
rect 64698 148294 64768 148350
rect 64448 148226 64768 148294
rect 64448 148170 64518 148226
rect 64574 148170 64642 148226
rect 64698 148170 64768 148226
rect 64448 148102 64768 148170
rect 64448 148046 64518 148102
rect 64574 148046 64642 148102
rect 64698 148046 64768 148102
rect 64448 147978 64768 148046
rect 64448 147922 64518 147978
rect 64574 147922 64642 147978
rect 64698 147922 64768 147978
rect 64448 147888 64768 147922
rect 95168 148350 95488 148384
rect 95168 148294 95238 148350
rect 95294 148294 95362 148350
rect 95418 148294 95488 148350
rect 95168 148226 95488 148294
rect 95168 148170 95238 148226
rect 95294 148170 95362 148226
rect 95418 148170 95488 148226
rect 95168 148102 95488 148170
rect 95168 148046 95238 148102
rect 95294 148046 95362 148102
rect 95418 148046 95488 148102
rect 95168 147978 95488 148046
rect 95168 147922 95238 147978
rect 95294 147922 95362 147978
rect 95418 147922 95488 147978
rect 95168 147888 95488 147922
rect 125888 148350 126208 148384
rect 125888 148294 125958 148350
rect 126014 148294 126082 148350
rect 126138 148294 126208 148350
rect 125888 148226 126208 148294
rect 125888 148170 125958 148226
rect 126014 148170 126082 148226
rect 126138 148170 126208 148226
rect 125888 148102 126208 148170
rect 125888 148046 125958 148102
rect 126014 148046 126082 148102
rect 126138 148046 126208 148102
rect 125888 147978 126208 148046
rect 125888 147922 125958 147978
rect 126014 147922 126082 147978
rect 126138 147922 126208 147978
rect 125888 147888 126208 147922
rect 156608 148350 156928 148384
rect 156608 148294 156678 148350
rect 156734 148294 156802 148350
rect 156858 148294 156928 148350
rect 156608 148226 156928 148294
rect 156608 148170 156678 148226
rect 156734 148170 156802 148226
rect 156858 148170 156928 148226
rect 156608 148102 156928 148170
rect 156608 148046 156678 148102
rect 156734 148046 156802 148102
rect 156858 148046 156928 148102
rect 156608 147978 156928 148046
rect 156608 147922 156678 147978
rect 156734 147922 156802 147978
rect 156858 147922 156928 147978
rect 156608 147888 156928 147922
rect 187328 148350 187648 148384
rect 187328 148294 187398 148350
rect 187454 148294 187522 148350
rect 187578 148294 187648 148350
rect 187328 148226 187648 148294
rect 187328 148170 187398 148226
rect 187454 148170 187522 148226
rect 187578 148170 187648 148226
rect 187328 148102 187648 148170
rect 187328 148046 187398 148102
rect 187454 148046 187522 148102
rect 187578 148046 187648 148102
rect 187328 147978 187648 148046
rect 187328 147922 187398 147978
rect 187454 147922 187522 147978
rect 187578 147922 187648 147978
rect 187328 147888 187648 147922
rect 218048 148350 218368 148384
rect 218048 148294 218118 148350
rect 218174 148294 218242 148350
rect 218298 148294 218368 148350
rect 218048 148226 218368 148294
rect 218048 148170 218118 148226
rect 218174 148170 218242 148226
rect 218298 148170 218368 148226
rect 218048 148102 218368 148170
rect 218048 148046 218118 148102
rect 218174 148046 218242 148102
rect 218298 148046 218368 148102
rect 218048 147978 218368 148046
rect 218048 147922 218118 147978
rect 218174 147922 218242 147978
rect 218298 147922 218368 147978
rect 218048 147888 218368 147922
rect 248768 148350 249088 148384
rect 248768 148294 248838 148350
rect 248894 148294 248962 148350
rect 249018 148294 249088 148350
rect 248768 148226 249088 148294
rect 248768 148170 248838 148226
rect 248894 148170 248962 148226
rect 249018 148170 249088 148226
rect 248768 148102 249088 148170
rect 248768 148046 248838 148102
rect 248894 148046 248962 148102
rect 249018 148046 249088 148102
rect 248768 147978 249088 148046
rect 248768 147922 248838 147978
rect 248894 147922 248962 147978
rect 249018 147922 249088 147978
rect 248768 147888 249088 147922
rect 279488 148350 279808 148384
rect 279488 148294 279558 148350
rect 279614 148294 279682 148350
rect 279738 148294 279808 148350
rect 279488 148226 279808 148294
rect 279488 148170 279558 148226
rect 279614 148170 279682 148226
rect 279738 148170 279808 148226
rect 279488 148102 279808 148170
rect 279488 148046 279558 148102
rect 279614 148046 279682 148102
rect 279738 148046 279808 148102
rect 279488 147978 279808 148046
rect 279488 147922 279558 147978
rect 279614 147922 279682 147978
rect 279738 147922 279808 147978
rect 279488 147888 279808 147922
rect 310208 148350 310528 148384
rect 310208 148294 310278 148350
rect 310334 148294 310402 148350
rect 310458 148294 310528 148350
rect 310208 148226 310528 148294
rect 310208 148170 310278 148226
rect 310334 148170 310402 148226
rect 310458 148170 310528 148226
rect 310208 148102 310528 148170
rect 310208 148046 310278 148102
rect 310334 148046 310402 148102
rect 310458 148046 310528 148102
rect 310208 147978 310528 148046
rect 310208 147922 310278 147978
rect 310334 147922 310402 147978
rect 310458 147922 310528 147978
rect 310208 147888 310528 147922
rect 340928 148350 341248 148384
rect 340928 148294 340998 148350
rect 341054 148294 341122 148350
rect 341178 148294 341248 148350
rect 340928 148226 341248 148294
rect 340928 148170 340998 148226
rect 341054 148170 341122 148226
rect 341178 148170 341248 148226
rect 340928 148102 341248 148170
rect 340928 148046 340998 148102
rect 341054 148046 341122 148102
rect 341178 148046 341248 148102
rect 340928 147978 341248 148046
rect 340928 147922 340998 147978
rect 341054 147922 341122 147978
rect 341178 147922 341248 147978
rect 340928 147888 341248 147922
rect 79808 136350 80128 136384
rect 79808 136294 79878 136350
rect 79934 136294 80002 136350
rect 80058 136294 80128 136350
rect 79808 136226 80128 136294
rect 79808 136170 79878 136226
rect 79934 136170 80002 136226
rect 80058 136170 80128 136226
rect 79808 136102 80128 136170
rect 79808 136046 79878 136102
rect 79934 136046 80002 136102
rect 80058 136046 80128 136102
rect 79808 135978 80128 136046
rect 79808 135922 79878 135978
rect 79934 135922 80002 135978
rect 80058 135922 80128 135978
rect 79808 135888 80128 135922
rect 110528 136350 110848 136384
rect 110528 136294 110598 136350
rect 110654 136294 110722 136350
rect 110778 136294 110848 136350
rect 110528 136226 110848 136294
rect 110528 136170 110598 136226
rect 110654 136170 110722 136226
rect 110778 136170 110848 136226
rect 110528 136102 110848 136170
rect 110528 136046 110598 136102
rect 110654 136046 110722 136102
rect 110778 136046 110848 136102
rect 110528 135978 110848 136046
rect 110528 135922 110598 135978
rect 110654 135922 110722 135978
rect 110778 135922 110848 135978
rect 110528 135888 110848 135922
rect 141248 136350 141568 136384
rect 141248 136294 141318 136350
rect 141374 136294 141442 136350
rect 141498 136294 141568 136350
rect 141248 136226 141568 136294
rect 141248 136170 141318 136226
rect 141374 136170 141442 136226
rect 141498 136170 141568 136226
rect 141248 136102 141568 136170
rect 141248 136046 141318 136102
rect 141374 136046 141442 136102
rect 141498 136046 141568 136102
rect 141248 135978 141568 136046
rect 141248 135922 141318 135978
rect 141374 135922 141442 135978
rect 141498 135922 141568 135978
rect 141248 135888 141568 135922
rect 171968 136350 172288 136384
rect 171968 136294 172038 136350
rect 172094 136294 172162 136350
rect 172218 136294 172288 136350
rect 171968 136226 172288 136294
rect 171968 136170 172038 136226
rect 172094 136170 172162 136226
rect 172218 136170 172288 136226
rect 171968 136102 172288 136170
rect 171968 136046 172038 136102
rect 172094 136046 172162 136102
rect 172218 136046 172288 136102
rect 171968 135978 172288 136046
rect 171968 135922 172038 135978
rect 172094 135922 172162 135978
rect 172218 135922 172288 135978
rect 171968 135888 172288 135922
rect 202688 136350 203008 136384
rect 202688 136294 202758 136350
rect 202814 136294 202882 136350
rect 202938 136294 203008 136350
rect 202688 136226 203008 136294
rect 202688 136170 202758 136226
rect 202814 136170 202882 136226
rect 202938 136170 203008 136226
rect 202688 136102 203008 136170
rect 202688 136046 202758 136102
rect 202814 136046 202882 136102
rect 202938 136046 203008 136102
rect 202688 135978 203008 136046
rect 202688 135922 202758 135978
rect 202814 135922 202882 135978
rect 202938 135922 203008 135978
rect 202688 135888 203008 135922
rect 233408 136350 233728 136384
rect 233408 136294 233478 136350
rect 233534 136294 233602 136350
rect 233658 136294 233728 136350
rect 233408 136226 233728 136294
rect 233408 136170 233478 136226
rect 233534 136170 233602 136226
rect 233658 136170 233728 136226
rect 233408 136102 233728 136170
rect 233408 136046 233478 136102
rect 233534 136046 233602 136102
rect 233658 136046 233728 136102
rect 233408 135978 233728 136046
rect 233408 135922 233478 135978
rect 233534 135922 233602 135978
rect 233658 135922 233728 135978
rect 233408 135888 233728 135922
rect 264128 136350 264448 136384
rect 264128 136294 264198 136350
rect 264254 136294 264322 136350
rect 264378 136294 264448 136350
rect 264128 136226 264448 136294
rect 264128 136170 264198 136226
rect 264254 136170 264322 136226
rect 264378 136170 264448 136226
rect 264128 136102 264448 136170
rect 264128 136046 264198 136102
rect 264254 136046 264322 136102
rect 264378 136046 264448 136102
rect 264128 135978 264448 136046
rect 264128 135922 264198 135978
rect 264254 135922 264322 135978
rect 264378 135922 264448 135978
rect 264128 135888 264448 135922
rect 294848 136350 295168 136384
rect 294848 136294 294918 136350
rect 294974 136294 295042 136350
rect 295098 136294 295168 136350
rect 294848 136226 295168 136294
rect 294848 136170 294918 136226
rect 294974 136170 295042 136226
rect 295098 136170 295168 136226
rect 294848 136102 295168 136170
rect 294848 136046 294918 136102
rect 294974 136046 295042 136102
rect 295098 136046 295168 136102
rect 294848 135978 295168 136046
rect 294848 135922 294918 135978
rect 294974 135922 295042 135978
rect 295098 135922 295168 135978
rect 294848 135888 295168 135922
rect 325568 136350 325888 136384
rect 325568 136294 325638 136350
rect 325694 136294 325762 136350
rect 325818 136294 325888 136350
rect 325568 136226 325888 136294
rect 325568 136170 325638 136226
rect 325694 136170 325762 136226
rect 325818 136170 325888 136226
rect 325568 136102 325888 136170
rect 325568 136046 325638 136102
rect 325694 136046 325762 136102
rect 325818 136046 325888 136102
rect 325568 135978 325888 136046
rect 325568 135922 325638 135978
rect 325694 135922 325762 135978
rect 325818 135922 325888 135978
rect 325568 135888 325888 135922
rect 348874 136350 349494 153922
rect 356288 154350 356608 154384
rect 356288 154294 356358 154350
rect 356414 154294 356482 154350
rect 356538 154294 356608 154350
rect 356288 154226 356608 154294
rect 356288 154170 356358 154226
rect 356414 154170 356482 154226
rect 356538 154170 356608 154226
rect 356288 154102 356608 154170
rect 356288 154046 356358 154102
rect 356414 154046 356482 154102
rect 356538 154046 356608 154102
rect 356288 153978 356608 154046
rect 356288 153922 356358 153978
rect 356414 153922 356482 153978
rect 356538 153922 356608 153978
rect 356288 153888 356608 153922
rect 363154 148350 363774 165922
rect 363154 148294 363250 148350
rect 363306 148294 363374 148350
rect 363430 148294 363498 148350
rect 363554 148294 363622 148350
rect 363678 148294 363774 148350
rect 363154 148226 363774 148294
rect 363154 148170 363250 148226
rect 363306 148170 363374 148226
rect 363430 148170 363498 148226
rect 363554 148170 363622 148226
rect 363678 148170 363774 148226
rect 363154 148102 363774 148170
rect 363154 148046 363250 148102
rect 363306 148046 363374 148102
rect 363430 148046 363498 148102
rect 363554 148046 363622 148102
rect 363678 148046 363774 148102
rect 363154 147978 363774 148046
rect 363154 147922 363250 147978
rect 363306 147922 363374 147978
rect 363430 147922 363498 147978
rect 363554 147922 363622 147978
rect 363678 147922 363774 147978
rect 348874 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 349494 136350
rect 348874 136226 349494 136294
rect 348874 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 349494 136226
rect 348874 136102 349494 136170
rect 348874 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 349494 136102
rect 348874 135978 349494 136046
rect 348874 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 349494 135978
rect 57154 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 57774 130350
rect 57154 130226 57774 130294
rect 57154 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 57774 130226
rect 57154 130102 57774 130170
rect 57154 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 57774 130102
rect 57154 129978 57774 130046
rect 57154 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 57774 129978
rect 57154 112350 57774 129922
rect 64448 130350 64768 130384
rect 64448 130294 64518 130350
rect 64574 130294 64642 130350
rect 64698 130294 64768 130350
rect 64448 130226 64768 130294
rect 64448 130170 64518 130226
rect 64574 130170 64642 130226
rect 64698 130170 64768 130226
rect 64448 130102 64768 130170
rect 64448 130046 64518 130102
rect 64574 130046 64642 130102
rect 64698 130046 64768 130102
rect 64448 129978 64768 130046
rect 64448 129922 64518 129978
rect 64574 129922 64642 129978
rect 64698 129922 64768 129978
rect 64448 129888 64768 129922
rect 95168 130350 95488 130384
rect 95168 130294 95238 130350
rect 95294 130294 95362 130350
rect 95418 130294 95488 130350
rect 95168 130226 95488 130294
rect 95168 130170 95238 130226
rect 95294 130170 95362 130226
rect 95418 130170 95488 130226
rect 95168 130102 95488 130170
rect 95168 130046 95238 130102
rect 95294 130046 95362 130102
rect 95418 130046 95488 130102
rect 95168 129978 95488 130046
rect 95168 129922 95238 129978
rect 95294 129922 95362 129978
rect 95418 129922 95488 129978
rect 95168 129888 95488 129922
rect 125888 130350 126208 130384
rect 125888 130294 125958 130350
rect 126014 130294 126082 130350
rect 126138 130294 126208 130350
rect 125888 130226 126208 130294
rect 125888 130170 125958 130226
rect 126014 130170 126082 130226
rect 126138 130170 126208 130226
rect 125888 130102 126208 130170
rect 125888 130046 125958 130102
rect 126014 130046 126082 130102
rect 126138 130046 126208 130102
rect 125888 129978 126208 130046
rect 125888 129922 125958 129978
rect 126014 129922 126082 129978
rect 126138 129922 126208 129978
rect 125888 129888 126208 129922
rect 156608 130350 156928 130384
rect 156608 130294 156678 130350
rect 156734 130294 156802 130350
rect 156858 130294 156928 130350
rect 156608 130226 156928 130294
rect 156608 130170 156678 130226
rect 156734 130170 156802 130226
rect 156858 130170 156928 130226
rect 156608 130102 156928 130170
rect 156608 130046 156678 130102
rect 156734 130046 156802 130102
rect 156858 130046 156928 130102
rect 156608 129978 156928 130046
rect 156608 129922 156678 129978
rect 156734 129922 156802 129978
rect 156858 129922 156928 129978
rect 156608 129888 156928 129922
rect 187328 130350 187648 130384
rect 187328 130294 187398 130350
rect 187454 130294 187522 130350
rect 187578 130294 187648 130350
rect 187328 130226 187648 130294
rect 187328 130170 187398 130226
rect 187454 130170 187522 130226
rect 187578 130170 187648 130226
rect 187328 130102 187648 130170
rect 187328 130046 187398 130102
rect 187454 130046 187522 130102
rect 187578 130046 187648 130102
rect 187328 129978 187648 130046
rect 187328 129922 187398 129978
rect 187454 129922 187522 129978
rect 187578 129922 187648 129978
rect 187328 129888 187648 129922
rect 218048 130350 218368 130384
rect 218048 130294 218118 130350
rect 218174 130294 218242 130350
rect 218298 130294 218368 130350
rect 218048 130226 218368 130294
rect 218048 130170 218118 130226
rect 218174 130170 218242 130226
rect 218298 130170 218368 130226
rect 218048 130102 218368 130170
rect 218048 130046 218118 130102
rect 218174 130046 218242 130102
rect 218298 130046 218368 130102
rect 218048 129978 218368 130046
rect 218048 129922 218118 129978
rect 218174 129922 218242 129978
rect 218298 129922 218368 129978
rect 218048 129888 218368 129922
rect 248768 130350 249088 130384
rect 248768 130294 248838 130350
rect 248894 130294 248962 130350
rect 249018 130294 249088 130350
rect 248768 130226 249088 130294
rect 248768 130170 248838 130226
rect 248894 130170 248962 130226
rect 249018 130170 249088 130226
rect 248768 130102 249088 130170
rect 248768 130046 248838 130102
rect 248894 130046 248962 130102
rect 249018 130046 249088 130102
rect 248768 129978 249088 130046
rect 248768 129922 248838 129978
rect 248894 129922 248962 129978
rect 249018 129922 249088 129978
rect 248768 129888 249088 129922
rect 279488 130350 279808 130384
rect 279488 130294 279558 130350
rect 279614 130294 279682 130350
rect 279738 130294 279808 130350
rect 279488 130226 279808 130294
rect 279488 130170 279558 130226
rect 279614 130170 279682 130226
rect 279738 130170 279808 130226
rect 279488 130102 279808 130170
rect 279488 130046 279558 130102
rect 279614 130046 279682 130102
rect 279738 130046 279808 130102
rect 279488 129978 279808 130046
rect 279488 129922 279558 129978
rect 279614 129922 279682 129978
rect 279738 129922 279808 129978
rect 279488 129888 279808 129922
rect 310208 130350 310528 130384
rect 310208 130294 310278 130350
rect 310334 130294 310402 130350
rect 310458 130294 310528 130350
rect 310208 130226 310528 130294
rect 310208 130170 310278 130226
rect 310334 130170 310402 130226
rect 310458 130170 310528 130226
rect 310208 130102 310528 130170
rect 310208 130046 310278 130102
rect 310334 130046 310402 130102
rect 310458 130046 310528 130102
rect 310208 129978 310528 130046
rect 310208 129922 310278 129978
rect 310334 129922 310402 129978
rect 310458 129922 310528 129978
rect 310208 129888 310528 129922
rect 340928 130350 341248 130384
rect 340928 130294 340998 130350
rect 341054 130294 341122 130350
rect 341178 130294 341248 130350
rect 340928 130226 341248 130294
rect 340928 130170 340998 130226
rect 341054 130170 341122 130226
rect 341178 130170 341248 130226
rect 340928 130102 341248 130170
rect 340928 130046 340998 130102
rect 341054 130046 341122 130102
rect 341178 130046 341248 130102
rect 340928 129978 341248 130046
rect 340928 129922 340998 129978
rect 341054 129922 341122 129978
rect 341178 129922 341248 129978
rect 340928 129888 341248 129922
rect 79808 118350 80128 118384
rect 79808 118294 79878 118350
rect 79934 118294 80002 118350
rect 80058 118294 80128 118350
rect 79808 118226 80128 118294
rect 79808 118170 79878 118226
rect 79934 118170 80002 118226
rect 80058 118170 80128 118226
rect 79808 118102 80128 118170
rect 79808 118046 79878 118102
rect 79934 118046 80002 118102
rect 80058 118046 80128 118102
rect 79808 117978 80128 118046
rect 79808 117922 79878 117978
rect 79934 117922 80002 117978
rect 80058 117922 80128 117978
rect 79808 117888 80128 117922
rect 110528 118350 110848 118384
rect 110528 118294 110598 118350
rect 110654 118294 110722 118350
rect 110778 118294 110848 118350
rect 110528 118226 110848 118294
rect 110528 118170 110598 118226
rect 110654 118170 110722 118226
rect 110778 118170 110848 118226
rect 110528 118102 110848 118170
rect 110528 118046 110598 118102
rect 110654 118046 110722 118102
rect 110778 118046 110848 118102
rect 110528 117978 110848 118046
rect 110528 117922 110598 117978
rect 110654 117922 110722 117978
rect 110778 117922 110848 117978
rect 110528 117888 110848 117922
rect 141248 118350 141568 118384
rect 141248 118294 141318 118350
rect 141374 118294 141442 118350
rect 141498 118294 141568 118350
rect 141248 118226 141568 118294
rect 141248 118170 141318 118226
rect 141374 118170 141442 118226
rect 141498 118170 141568 118226
rect 141248 118102 141568 118170
rect 141248 118046 141318 118102
rect 141374 118046 141442 118102
rect 141498 118046 141568 118102
rect 141248 117978 141568 118046
rect 141248 117922 141318 117978
rect 141374 117922 141442 117978
rect 141498 117922 141568 117978
rect 141248 117888 141568 117922
rect 171968 118350 172288 118384
rect 171968 118294 172038 118350
rect 172094 118294 172162 118350
rect 172218 118294 172288 118350
rect 171968 118226 172288 118294
rect 171968 118170 172038 118226
rect 172094 118170 172162 118226
rect 172218 118170 172288 118226
rect 171968 118102 172288 118170
rect 171968 118046 172038 118102
rect 172094 118046 172162 118102
rect 172218 118046 172288 118102
rect 171968 117978 172288 118046
rect 171968 117922 172038 117978
rect 172094 117922 172162 117978
rect 172218 117922 172288 117978
rect 171968 117888 172288 117922
rect 202688 118350 203008 118384
rect 202688 118294 202758 118350
rect 202814 118294 202882 118350
rect 202938 118294 203008 118350
rect 202688 118226 203008 118294
rect 202688 118170 202758 118226
rect 202814 118170 202882 118226
rect 202938 118170 203008 118226
rect 202688 118102 203008 118170
rect 202688 118046 202758 118102
rect 202814 118046 202882 118102
rect 202938 118046 203008 118102
rect 202688 117978 203008 118046
rect 202688 117922 202758 117978
rect 202814 117922 202882 117978
rect 202938 117922 203008 117978
rect 202688 117888 203008 117922
rect 233408 118350 233728 118384
rect 233408 118294 233478 118350
rect 233534 118294 233602 118350
rect 233658 118294 233728 118350
rect 233408 118226 233728 118294
rect 233408 118170 233478 118226
rect 233534 118170 233602 118226
rect 233658 118170 233728 118226
rect 233408 118102 233728 118170
rect 233408 118046 233478 118102
rect 233534 118046 233602 118102
rect 233658 118046 233728 118102
rect 233408 117978 233728 118046
rect 233408 117922 233478 117978
rect 233534 117922 233602 117978
rect 233658 117922 233728 117978
rect 233408 117888 233728 117922
rect 264128 118350 264448 118384
rect 264128 118294 264198 118350
rect 264254 118294 264322 118350
rect 264378 118294 264448 118350
rect 264128 118226 264448 118294
rect 264128 118170 264198 118226
rect 264254 118170 264322 118226
rect 264378 118170 264448 118226
rect 264128 118102 264448 118170
rect 264128 118046 264198 118102
rect 264254 118046 264322 118102
rect 264378 118046 264448 118102
rect 264128 117978 264448 118046
rect 264128 117922 264198 117978
rect 264254 117922 264322 117978
rect 264378 117922 264448 117978
rect 264128 117888 264448 117922
rect 294848 118350 295168 118384
rect 294848 118294 294918 118350
rect 294974 118294 295042 118350
rect 295098 118294 295168 118350
rect 294848 118226 295168 118294
rect 294848 118170 294918 118226
rect 294974 118170 295042 118226
rect 295098 118170 295168 118226
rect 294848 118102 295168 118170
rect 294848 118046 294918 118102
rect 294974 118046 295042 118102
rect 295098 118046 295168 118102
rect 294848 117978 295168 118046
rect 294848 117922 294918 117978
rect 294974 117922 295042 117978
rect 295098 117922 295168 117978
rect 294848 117888 295168 117922
rect 325568 118350 325888 118384
rect 325568 118294 325638 118350
rect 325694 118294 325762 118350
rect 325818 118294 325888 118350
rect 325568 118226 325888 118294
rect 325568 118170 325638 118226
rect 325694 118170 325762 118226
rect 325818 118170 325888 118226
rect 325568 118102 325888 118170
rect 325568 118046 325638 118102
rect 325694 118046 325762 118102
rect 325818 118046 325888 118102
rect 325568 117978 325888 118046
rect 325568 117922 325638 117978
rect 325694 117922 325762 117978
rect 325818 117922 325888 117978
rect 325568 117888 325888 117922
rect 348874 118350 349494 135922
rect 356288 136350 356608 136384
rect 356288 136294 356358 136350
rect 356414 136294 356482 136350
rect 356538 136294 356608 136350
rect 356288 136226 356608 136294
rect 356288 136170 356358 136226
rect 356414 136170 356482 136226
rect 356538 136170 356608 136226
rect 356288 136102 356608 136170
rect 356288 136046 356358 136102
rect 356414 136046 356482 136102
rect 356538 136046 356608 136102
rect 356288 135978 356608 136046
rect 356288 135922 356358 135978
rect 356414 135922 356482 135978
rect 356538 135922 356608 135978
rect 356288 135888 356608 135922
rect 363154 130350 363774 147922
rect 363154 130294 363250 130350
rect 363306 130294 363374 130350
rect 363430 130294 363498 130350
rect 363554 130294 363622 130350
rect 363678 130294 363774 130350
rect 363154 130226 363774 130294
rect 363154 130170 363250 130226
rect 363306 130170 363374 130226
rect 363430 130170 363498 130226
rect 363554 130170 363622 130226
rect 363678 130170 363774 130226
rect 363154 130102 363774 130170
rect 363154 130046 363250 130102
rect 363306 130046 363374 130102
rect 363430 130046 363498 130102
rect 363554 130046 363622 130102
rect 363678 130046 363774 130102
rect 363154 129978 363774 130046
rect 363154 129922 363250 129978
rect 363306 129922 363374 129978
rect 363430 129922 363498 129978
rect 363554 129922 363622 129978
rect 363678 129922 363774 129978
rect 348874 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 349494 118350
rect 348874 118226 349494 118294
rect 348874 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 349494 118226
rect 348874 118102 349494 118170
rect 348874 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 349494 118102
rect 348874 117978 349494 118046
rect 348874 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 349494 117978
rect 57154 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 57774 112350
rect 57154 112226 57774 112294
rect 57154 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 57774 112226
rect 57154 112102 57774 112170
rect 57154 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 57774 112102
rect 57154 111978 57774 112046
rect 57154 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 57774 111978
rect 57154 94350 57774 111922
rect 64448 112350 64768 112384
rect 64448 112294 64518 112350
rect 64574 112294 64642 112350
rect 64698 112294 64768 112350
rect 64448 112226 64768 112294
rect 64448 112170 64518 112226
rect 64574 112170 64642 112226
rect 64698 112170 64768 112226
rect 64448 112102 64768 112170
rect 64448 112046 64518 112102
rect 64574 112046 64642 112102
rect 64698 112046 64768 112102
rect 64448 111978 64768 112046
rect 64448 111922 64518 111978
rect 64574 111922 64642 111978
rect 64698 111922 64768 111978
rect 64448 111888 64768 111922
rect 95168 112350 95488 112384
rect 95168 112294 95238 112350
rect 95294 112294 95362 112350
rect 95418 112294 95488 112350
rect 95168 112226 95488 112294
rect 95168 112170 95238 112226
rect 95294 112170 95362 112226
rect 95418 112170 95488 112226
rect 95168 112102 95488 112170
rect 95168 112046 95238 112102
rect 95294 112046 95362 112102
rect 95418 112046 95488 112102
rect 95168 111978 95488 112046
rect 95168 111922 95238 111978
rect 95294 111922 95362 111978
rect 95418 111922 95488 111978
rect 95168 111888 95488 111922
rect 125888 112350 126208 112384
rect 125888 112294 125958 112350
rect 126014 112294 126082 112350
rect 126138 112294 126208 112350
rect 125888 112226 126208 112294
rect 125888 112170 125958 112226
rect 126014 112170 126082 112226
rect 126138 112170 126208 112226
rect 125888 112102 126208 112170
rect 125888 112046 125958 112102
rect 126014 112046 126082 112102
rect 126138 112046 126208 112102
rect 125888 111978 126208 112046
rect 125888 111922 125958 111978
rect 126014 111922 126082 111978
rect 126138 111922 126208 111978
rect 125888 111888 126208 111922
rect 156608 112350 156928 112384
rect 156608 112294 156678 112350
rect 156734 112294 156802 112350
rect 156858 112294 156928 112350
rect 156608 112226 156928 112294
rect 156608 112170 156678 112226
rect 156734 112170 156802 112226
rect 156858 112170 156928 112226
rect 156608 112102 156928 112170
rect 156608 112046 156678 112102
rect 156734 112046 156802 112102
rect 156858 112046 156928 112102
rect 156608 111978 156928 112046
rect 156608 111922 156678 111978
rect 156734 111922 156802 111978
rect 156858 111922 156928 111978
rect 156608 111888 156928 111922
rect 187328 112350 187648 112384
rect 187328 112294 187398 112350
rect 187454 112294 187522 112350
rect 187578 112294 187648 112350
rect 187328 112226 187648 112294
rect 187328 112170 187398 112226
rect 187454 112170 187522 112226
rect 187578 112170 187648 112226
rect 187328 112102 187648 112170
rect 187328 112046 187398 112102
rect 187454 112046 187522 112102
rect 187578 112046 187648 112102
rect 187328 111978 187648 112046
rect 187328 111922 187398 111978
rect 187454 111922 187522 111978
rect 187578 111922 187648 111978
rect 187328 111888 187648 111922
rect 218048 112350 218368 112384
rect 218048 112294 218118 112350
rect 218174 112294 218242 112350
rect 218298 112294 218368 112350
rect 218048 112226 218368 112294
rect 218048 112170 218118 112226
rect 218174 112170 218242 112226
rect 218298 112170 218368 112226
rect 218048 112102 218368 112170
rect 218048 112046 218118 112102
rect 218174 112046 218242 112102
rect 218298 112046 218368 112102
rect 218048 111978 218368 112046
rect 218048 111922 218118 111978
rect 218174 111922 218242 111978
rect 218298 111922 218368 111978
rect 218048 111888 218368 111922
rect 248768 112350 249088 112384
rect 248768 112294 248838 112350
rect 248894 112294 248962 112350
rect 249018 112294 249088 112350
rect 248768 112226 249088 112294
rect 248768 112170 248838 112226
rect 248894 112170 248962 112226
rect 249018 112170 249088 112226
rect 248768 112102 249088 112170
rect 248768 112046 248838 112102
rect 248894 112046 248962 112102
rect 249018 112046 249088 112102
rect 248768 111978 249088 112046
rect 248768 111922 248838 111978
rect 248894 111922 248962 111978
rect 249018 111922 249088 111978
rect 248768 111888 249088 111922
rect 279488 112350 279808 112384
rect 279488 112294 279558 112350
rect 279614 112294 279682 112350
rect 279738 112294 279808 112350
rect 279488 112226 279808 112294
rect 279488 112170 279558 112226
rect 279614 112170 279682 112226
rect 279738 112170 279808 112226
rect 279488 112102 279808 112170
rect 279488 112046 279558 112102
rect 279614 112046 279682 112102
rect 279738 112046 279808 112102
rect 279488 111978 279808 112046
rect 279488 111922 279558 111978
rect 279614 111922 279682 111978
rect 279738 111922 279808 111978
rect 279488 111888 279808 111922
rect 310208 112350 310528 112384
rect 310208 112294 310278 112350
rect 310334 112294 310402 112350
rect 310458 112294 310528 112350
rect 310208 112226 310528 112294
rect 310208 112170 310278 112226
rect 310334 112170 310402 112226
rect 310458 112170 310528 112226
rect 310208 112102 310528 112170
rect 310208 112046 310278 112102
rect 310334 112046 310402 112102
rect 310458 112046 310528 112102
rect 310208 111978 310528 112046
rect 310208 111922 310278 111978
rect 310334 111922 310402 111978
rect 310458 111922 310528 111978
rect 310208 111888 310528 111922
rect 340928 112350 341248 112384
rect 340928 112294 340998 112350
rect 341054 112294 341122 112350
rect 341178 112294 341248 112350
rect 340928 112226 341248 112294
rect 340928 112170 340998 112226
rect 341054 112170 341122 112226
rect 341178 112170 341248 112226
rect 340928 112102 341248 112170
rect 340928 112046 340998 112102
rect 341054 112046 341122 112102
rect 341178 112046 341248 112102
rect 340928 111978 341248 112046
rect 340928 111922 340998 111978
rect 341054 111922 341122 111978
rect 341178 111922 341248 111978
rect 340928 111888 341248 111922
rect 79808 100350 80128 100384
rect 79808 100294 79878 100350
rect 79934 100294 80002 100350
rect 80058 100294 80128 100350
rect 79808 100226 80128 100294
rect 79808 100170 79878 100226
rect 79934 100170 80002 100226
rect 80058 100170 80128 100226
rect 79808 100102 80128 100170
rect 79808 100046 79878 100102
rect 79934 100046 80002 100102
rect 80058 100046 80128 100102
rect 79808 99978 80128 100046
rect 79808 99922 79878 99978
rect 79934 99922 80002 99978
rect 80058 99922 80128 99978
rect 79808 99888 80128 99922
rect 110528 100350 110848 100384
rect 110528 100294 110598 100350
rect 110654 100294 110722 100350
rect 110778 100294 110848 100350
rect 110528 100226 110848 100294
rect 110528 100170 110598 100226
rect 110654 100170 110722 100226
rect 110778 100170 110848 100226
rect 110528 100102 110848 100170
rect 110528 100046 110598 100102
rect 110654 100046 110722 100102
rect 110778 100046 110848 100102
rect 110528 99978 110848 100046
rect 110528 99922 110598 99978
rect 110654 99922 110722 99978
rect 110778 99922 110848 99978
rect 110528 99888 110848 99922
rect 141248 100350 141568 100384
rect 141248 100294 141318 100350
rect 141374 100294 141442 100350
rect 141498 100294 141568 100350
rect 141248 100226 141568 100294
rect 141248 100170 141318 100226
rect 141374 100170 141442 100226
rect 141498 100170 141568 100226
rect 141248 100102 141568 100170
rect 141248 100046 141318 100102
rect 141374 100046 141442 100102
rect 141498 100046 141568 100102
rect 141248 99978 141568 100046
rect 141248 99922 141318 99978
rect 141374 99922 141442 99978
rect 141498 99922 141568 99978
rect 141248 99888 141568 99922
rect 171968 100350 172288 100384
rect 171968 100294 172038 100350
rect 172094 100294 172162 100350
rect 172218 100294 172288 100350
rect 171968 100226 172288 100294
rect 171968 100170 172038 100226
rect 172094 100170 172162 100226
rect 172218 100170 172288 100226
rect 171968 100102 172288 100170
rect 171968 100046 172038 100102
rect 172094 100046 172162 100102
rect 172218 100046 172288 100102
rect 171968 99978 172288 100046
rect 171968 99922 172038 99978
rect 172094 99922 172162 99978
rect 172218 99922 172288 99978
rect 171968 99888 172288 99922
rect 202688 100350 203008 100384
rect 202688 100294 202758 100350
rect 202814 100294 202882 100350
rect 202938 100294 203008 100350
rect 202688 100226 203008 100294
rect 202688 100170 202758 100226
rect 202814 100170 202882 100226
rect 202938 100170 203008 100226
rect 202688 100102 203008 100170
rect 202688 100046 202758 100102
rect 202814 100046 202882 100102
rect 202938 100046 203008 100102
rect 202688 99978 203008 100046
rect 202688 99922 202758 99978
rect 202814 99922 202882 99978
rect 202938 99922 203008 99978
rect 202688 99888 203008 99922
rect 233408 100350 233728 100384
rect 233408 100294 233478 100350
rect 233534 100294 233602 100350
rect 233658 100294 233728 100350
rect 233408 100226 233728 100294
rect 233408 100170 233478 100226
rect 233534 100170 233602 100226
rect 233658 100170 233728 100226
rect 233408 100102 233728 100170
rect 233408 100046 233478 100102
rect 233534 100046 233602 100102
rect 233658 100046 233728 100102
rect 233408 99978 233728 100046
rect 233408 99922 233478 99978
rect 233534 99922 233602 99978
rect 233658 99922 233728 99978
rect 233408 99888 233728 99922
rect 264128 100350 264448 100384
rect 264128 100294 264198 100350
rect 264254 100294 264322 100350
rect 264378 100294 264448 100350
rect 264128 100226 264448 100294
rect 264128 100170 264198 100226
rect 264254 100170 264322 100226
rect 264378 100170 264448 100226
rect 264128 100102 264448 100170
rect 264128 100046 264198 100102
rect 264254 100046 264322 100102
rect 264378 100046 264448 100102
rect 264128 99978 264448 100046
rect 264128 99922 264198 99978
rect 264254 99922 264322 99978
rect 264378 99922 264448 99978
rect 264128 99888 264448 99922
rect 294848 100350 295168 100384
rect 294848 100294 294918 100350
rect 294974 100294 295042 100350
rect 295098 100294 295168 100350
rect 294848 100226 295168 100294
rect 294848 100170 294918 100226
rect 294974 100170 295042 100226
rect 295098 100170 295168 100226
rect 294848 100102 295168 100170
rect 294848 100046 294918 100102
rect 294974 100046 295042 100102
rect 295098 100046 295168 100102
rect 294848 99978 295168 100046
rect 294848 99922 294918 99978
rect 294974 99922 295042 99978
rect 295098 99922 295168 99978
rect 294848 99888 295168 99922
rect 325568 100350 325888 100384
rect 325568 100294 325638 100350
rect 325694 100294 325762 100350
rect 325818 100294 325888 100350
rect 325568 100226 325888 100294
rect 325568 100170 325638 100226
rect 325694 100170 325762 100226
rect 325818 100170 325888 100226
rect 325568 100102 325888 100170
rect 325568 100046 325638 100102
rect 325694 100046 325762 100102
rect 325818 100046 325888 100102
rect 325568 99978 325888 100046
rect 325568 99922 325638 99978
rect 325694 99922 325762 99978
rect 325818 99922 325888 99978
rect 325568 99888 325888 99922
rect 348874 100350 349494 117922
rect 356288 118350 356608 118384
rect 356288 118294 356358 118350
rect 356414 118294 356482 118350
rect 356538 118294 356608 118350
rect 356288 118226 356608 118294
rect 356288 118170 356358 118226
rect 356414 118170 356482 118226
rect 356538 118170 356608 118226
rect 356288 118102 356608 118170
rect 356288 118046 356358 118102
rect 356414 118046 356482 118102
rect 356538 118046 356608 118102
rect 356288 117978 356608 118046
rect 356288 117922 356358 117978
rect 356414 117922 356482 117978
rect 356538 117922 356608 117978
rect 356288 117888 356608 117922
rect 363154 112350 363774 129922
rect 363154 112294 363250 112350
rect 363306 112294 363374 112350
rect 363430 112294 363498 112350
rect 363554 112294 363622 112350
rect 363678 112294 363774 112350
rect 363154 112226 363774 112294
rect 363154 112170 363250 112226
rect 363306 112170 363374 112226
rect 363430 112170 363498 112226
rect 363554 112170 363622 112226
rect 363678 112170 363774 112226
rect 363154 112102 363774 112170
rect 363154 112046 363250 112102
rect 363306 112046 363374 112102
rect 363430 112046 363498 112102
rect 363554 112046 363622 112102
rect 363678 112046 363774 112102
rect 363154 111978 363774 112046
rect 363154 111922 363250 111978
rect 363306 111922 363374 111978
rect 363430 111922 363498 111978
rect 363554 111922 363622 111978
rect 363678 111922 363774 111978
rect 348874 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 349494 100350
rect 348874 100226 349494 100294
rect 348874 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 349494 100226
rect 348874 100102 349494 100170
rect 348874 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 349494 100102
rect 348874 99978 349494 100046
rect 348874 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 349494 99978
rect 57154 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 57774 94350
rect 57154 94226 57774 94294
rect 57154 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 57774 94226
rect 57154 94102 57774 94170
rect 57154 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 57774 94102
rect 57154 93978 57774 94046
rect 57154 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 57774 93978
rect 57154 76350 57774 93922
rect 64448 94350 64768 94384
rect 64448 94294 64518 94350
rect 64574 94294 64642 94350
rect 64698 94294 64768 94350
rect 64448 94226 64768 94294
rect 64448 94170 64518 94226
rect 64574 94170 64642 94226
rect 64698 94170 64768 94226
rect 64448 94102 64768 94170
rect 64448 94046 64518 94102
rect 64574 94046 64642 94102
rect 64698 94046 64768 94102
rect 64448 93978 64768 94046
rect 64448 93922 64518 93978
rect 64574 93922 64642 93978
rect 64698 93922 64768 93978
rect 64448 93888 64768 93922
rect 95168 94350 95488 94384
rect 95168 94294 95238 94350
rect 95294 94294 95362 94350
rect 95418 94294 95488 94350
rect 95168 94226 95488 94294
rect 95168 94170 95238 94226
rect 95294 94170 95362 94226
rect 95418 94170 95488 94226
rect 95168 94102 95488 94170
rect 95168 94046 95238 94102
rect 95294 94046 95362 94102
rect 95418 94046 95488 94102
rect 95168 93978 95488 94046
rect 95168 93922 95238 93978
rect 95294 93922 95362 93978
rect 95418 93922 95488 93978
rect 95168 93888 95488 93922
rect 125888 94350 126208 94384
rect 125888 94294 125958 94350
rect 126014 94294 126082 94350
rect 126138 94294 126208 94350
rect 125888 94226 126208 94294
rect 125888 94170 125958 94226
rect 126014 94170 126082 94226
rect 126138 94170 126208 94226
rect 125888 94102 126208 94170
rect 125888 94046 125958 94102
rect 126014 94046 126082 94102
rect 126138 94046 126208 94102
rect 125888 93978 126208 94046
rect 125888 93922 125958 93978
rect 126014 93922 126082 93978
rect 126138 93922 126208 93978
rect 125888 93888 126208 93922
rect 156608 94350 156928 94384
rect 156608 94294 156678 94350
rect 156734 94294 156802 94350
rect 156858 94294 156928 94350
rect 156608 94226 156928 94294
rect 156608 94170 156678 94226
rect 156734 94170 156802 94226
rect 156858 94170 156928 94226
rect 156608 94102 156928 94170
rect 156608 94046 156678 94102
rect 156734 94046 156802 94102
rect 156858 94046 156928 94102
rect 156608 93978 156928 94046
rect 156608 93922 156678 93978
rect 156734 93922 156802 93978
rect 156858 93922 156928 93978
rect 156608 93888 156928 93922
rect 187328 94350 187648 94384
rect 187328 94294 187398 94350
rect 187454 94294 187522 94350
rect 187578 94294 187648 94350
rect 187328 94226 187648 94294
rect 187328 94170 187398 94226
rect 187454 94170 187522 94226
rect 187578 94170 187648 94226
rect 187328 94102 187648 94170
rect 187328 94046 187398 94102
rect 187454 94046 187522 94102
rect 187578 94046 187648 94102
rect 187328 93978 187648 94046
rect 187328 93922 187398 93978
rect 187454 93922 187522 93978
rect 187578 93922 187648 93978
rect 187328 93888 187648 93922
rect 218048 94350 218368 94384
rect 218048 94294 218118 94350
rect 218174 94294 218242 94350
rect 218298 94294 218368 94350
rect 218048 94226 218368 94294
rect 218048 94170 218118 94226
rect 218174 94170 218242 94226
rect 218298 94170 218368 94226
rect 218048 94102 218368 94170
rect 218048 94046 218118 94102
rect 218174 94046 218242 94102
rect 218298 94046 218368 94102
rect 218048 93978 218368 94046
rect 218048 93922 218118 93978
rect 218174 93922 218242 93978
rect 218298 93922 218368 93978
rect 218048 93888 218368 93922
rect 248768 94350 249088 94384
rect 248768 94294 248838 94350
rect 248894 94294 248962 94350
rect 249018 94294 249088 94350
rect 248768 94226 249088 94294
rect 248768 94170 248838 94226
rect 248894 94170 248962 94226
rect 249018 94170 249088 94226
rect 248768 94102 249088 94170
rect 248768 94046 248838 94102
rect 248894 94046 248962 94102
rect 249018 94046 249088 94102
rect 248768 93978 249088 94046
rect 248768 93922 248838 93978
rect 248894 93922 248962 93978
rect 249018 93922 249088 93978
rect 248768 93888 249088 93922
rect 279488 94350 279808 94384
rect 279488 94294 279558 94350
rect 279614 94294 279682 94350
rect 279738 94294 279808 94350
rect 279488 94226 279808 94294
rect 279488 94170 279558 94226
rect 279614 94170 279682 94226
rect 279738 94170 279808 94226
rect 279488 94102 279808 94170
rect 279488 94046 279558 94102
rect 279614 94046 279682 94102
rect 279738 94046 279808 94102
rect 279488 93978 279808 94046
rect 279488 93922 279558 93978
rect 279614 93922 279682 93978
rect 279738 93922 279808 93978
rect 279488 93888 279808 93922
rect 310208 94350 310528 94384
rect 310208 94294 310278 94350
rect 310334 94294 310402 94350
rect 310458 94294 310528 94350
rect 310208 94226 310528 94294
rect 310208 94170 310278 94226
rect 310334 94170 310402 94226
rect 310458 94170 310528 94226
rect 310208 94102 310528 94170
rect 310208 94046 310278 94102
rect 310334 94046 310402 94102
rect 310458 94046 310528 94102
rect 310208 93978 310528 94046
rect 310208 93922 310278 93978
rect 310334 93922 310402 93978
rect 310458 93922 310528 93978
rect 310208 93888 310528 93922
rect 340928 94350 341248 94384
rect 340928 94294 340998 94350
rect 341054 94294 341122 94350
rect 341178 94294 341248 94350
rect 340928 94226 341248 94294
rect 340928 94170 340998 94226
rect 341054 94170 341122 94226
rect 341178 94170 341248 94226
rect 340928 94102 341248 94170
rect 340928 94046 340998 94102
rect 341054 94046 341122 94102
rect 341178 94046 341248 94102
rect 340928 93978 341248 94046
rect 340928 93922 340998 93978
rect 341054 93922 341122 93978
rect 341178 93922 341248 93978
rect 340928 93888 341248 93922
rect 79808 82350 80128 82384
rect 79808 82294 79878 82350
rect 79934 82294 80002 82350
rect 80058 82294 80128 82350
rect 79808 82226 80128 82294
rect 79808 82170 79878 82226
rect 79934 82170 80002 82226
rect 80058 82170 80128 82226
rect 79808 82102 80128 82170
rect 79808 82046 79878 82102
rect 79934 82046 80002 82102
rect 80058 82046 80128 82102
rect 79808 81978 80128 82046
rect 79808 81922 79878 81978
rect 79934 81922 80002 81978
rect 80058 81922 80128 81978
rect 79808 81888 80128 81922
rect 110528 82350 110848 82384
rect 110528 82294 110598 82350
rect 110654 82294 110722 82350
rect 110778 82294 110848 82350
rect 110528 82226 110848 82294
rect 110528 82170 110598 82226
rect 110654 82170 110722 82226
rect 110778 82170 110848 82226
rect 110528 82102 110848 82170
rect 110528 82046 110598 82102
rect 110654 82046 110722 82102
rect 110778 82046 110848 82102
rect 110528 81978 110848 82046
rect 110528 81922 110598 81978
rect 110654 81922 110722 81978
rect 110778 81922 110848 81978
rect 110528 81888 110848 81922
rect 141248 82350 141568 82384
rect 141248 82294 141318 82350
rect 141374 82294 141442 82350
rect 141498 82294 141568 82350
rect 141248 82226 141568 82294
rect 141248 82170 141318 82226
rect 141374 82170 141442 82226
rect 141498 82170 141568 82226
rect 141248 82102 141568 82170
rect 141248 82046 141318 82102
rect 141374 82046 141442 82102
rect 141498 82046 141568 82102
rect 141248 81978 141568 82046
rect 141248 81922 141318 81978
rect 141374 81922 141442 81978
rect 141498 81922 141568 81978
rect 141248 81888 141568 81922
rect 171968 82350 172288 82384
rect 171968 82294 172038 82350
rect 172094 82294 172162 82350
rect 172218 82294 172288 82350
rect 171968 82226 172288 82294
rect 171968 82170 172038 82226
rect 172094 82170 172162 82226
rect 172218 82170 172288 82226
rect 171968 82102 172288 82170
rect 171968 82046 172038 82102
rect 172094 82046 172162 82102
rect 172218 82046 172288 82102
rect 171968 81978 172288 82046
rect 171968 81922 172038 81978
rect 172094 81922 172162 81978
rect 172218 81922 172288 81978
rect 171968 81888 172288 81922
rect 202688 82350 203008 82384
rect 202688 82294 202758 82350
rect 202814 82294 202882 82350
rect 202938 82294 203008 82350
rect 202688 82226 203008 82294
rect 202688 82170 202758 82226
rect 202814 82170 202882 82226
rect 202938 82170 203008 82226
rect 202688 82102 203008 82170
rect 202688 82046 202758 82102
rect 202814 82046 202882 82102
rect 202938 82046 203008 82102
rect 202688 81978 203008 82046
rect 202688 81922 202758 81978
rect 202814 81922 202882 81978
rect 202938 81922 203008 81978
rect 202688 81888 203008 81922
rect 233408 82350 233728 82384
rect 233408 82294 233478 82350
rect 233534 82294 233602 82350
rect 233658 82294 233728 82350
rect 233408 82226 233728 82294
rect 233408 82170 233478 82226
rect 233534 82170 233602 82226
rect 233658 82170 233728 82226
rect 233408 82102 233728 82170
rect 233408 82046 233478 82102
rect 233534 82046 233602 82102
rect 233658 82046 233728 82102
rect 233408 81978 233728 82046
rect 233408 81922 233478 81978
rect 233534 81922 233602 81978
rect 233658 81922 233728 81978
rect 233408 81888 233728 81922
rect 264128 82350 264448 82384
rect 264128 82294 264198 82350
rect 264254 82294 264322 82350
rect 264378 82294 264448 82350
rect 264128 82226 264448 82294
rect 264128 82170 264198 82226
rect 264254 82170 264322 82226
rect 264378 82170 264448 82226
rect 264128 82102 264448 82170
rect 264128 82046 264198 82102
rect 264254 82046 264322 82102
rect 264378 82046 264448 82102
rect 264128 81978 264448 82046
rect 264128 81922 264198 81978
rect 264254 81922 264322 81978
rect 264378 81922 264448 81978
rect 264128 81888 264448 81922
rect 294848 82350 295168 82384
rect 294848 82294 294918 82350
rect 294974 82294 295042 82350
rect 295098 82294 295168 82350
rect 294848 82226 295168 82294
rect 294848 82170 294918 82226
rect 294974 82170 295042 82226
rect 295098 82170 295168 82226
rect 294848 82102 295168 82170
rect 294848 82046 294918 82102
rect 294974 82046 295042 82102
rect 295098 82046 295168 82102
rect 294848 81978 295168 82046
rect 294848 81922 294918 81978
rect 294974 81922 295042 81978
rect 295098 81922 295168 81978
rect 294848 81888 295168 81922
rect 325568 82350 325888 82384
rect 325568 82294 325638 82350
rect 325694 82294 325762 82350
rect 325818 82294 325888 82350
rect 325568 82226 325888 82294
rect 325568 82170 325638 82226
rect 325694 82170 325762 82226
rect 325818 82170 325888 82226
rect 325568 82102 325888 82170
rect 325568 82046 325638 82102
rect 325694 82046 325762 82102
rect 325818 82046 325888 82102
rect 325568 81978 325888 82046
rect 325568 81922 325638 81978
rect 325694 81922 325762 81978
rect 325818 81922 325888 81978
rect 325568 81888 325888 81922
rect 348874 82350 349494 99922
rect 356288 100350 356608 100384
rect 356288 100294 356358 100350
rect 356414 100294 356482 100350
rect 356538 100294 356608 100350
rect 356288 100226 356608 100294
rect 356288 100170 356358 100226
rect 356414 100170 356482 100226
rect 356538 100170 356608 100226
rect 356288 100102 356608 100170
rect 356288 100046 356358 100102
rect 356414 100046 356482 100102
rect 356538 100046 356608 100102
rect 356288 99978 356608 100046
rect 356288 99922 356358 99978
rect 356414 99922 356482 99978
rect 356538 99922 356608 99978
rect 356288 99888 356608 99922
rect 363154 94350 363774 111922
rect 363154 94294 363250 94350
rect 363306 94294 363374 94350
rect 363430 94294 363498 94350
rect 363554 94294 363622 94350
rect 363678 94294 363774 94350
rect 363154 94226 363774 94294
rect 363154 94170 363250 94226
rect 363306 94170 363374 94226
rect 363430 94170 363498 94226
rect 363554 94170 363622 94226
rect 363678 94170 363774 94226
rect 363154 94102 363774 94170
rect 363154 94046 363250 94102
rect 363306 94046 363374 94102
rect 363430 94046 363498 94102
rect 363554 94046 363622 94102
rect 363678 94046 363774 94102
rect 363154 93978 363774 94046
rect 363154 93922 363250 93978
rect 363306 93922 363374 93978
rect 363430 93922 363498 93978
rect 363554 93922 363622 93978
rect 363678 93922 363774 93978
rect 348874 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 349494 82350
rect 348874 82226 349494 82294
rect 348874 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 349494 82226
rect 348874 82102 349494 82170
rect 348874 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 349494 82102
rect 348874 81978 349494 82046
rect 348874 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 349494 81978
rect 57154 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 57774 76350
rect 57154 76226 57774 76294
rect 57154 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 57774 76226
rect 57154 76102 57774 76170
rect 57154 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 57774 76102
rect 57154 75978 57774 76046
rect 57154 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 57774 75978
rect 57154 58350 57774 75922
rect 64448 76350 64768 76384
rect 64448 76294 64518 76350
rect 64574 76294 64642 76350
rect 64698 76294 64768 76350
rect 64448 76226 64768 76294
rect 64448 76170 64518 76226
rect 64574 76170 64642 76226
rect 64698 76170 64768 76226
rect 64448 76102 64768 76170
rect 64448 76046 64518 76102
rect 64574 76046 64642 76102
rect 64698 76046 64768 76102
rect 64448 75978 64768 76046
rect 64448 75922 64518 75978
rect 64574 75922 64642 75978
rect 64698 75922 64768 75978
rect 64448 75888 64768 75922
rect 95168 76350 95488 76384
rect 95168 76294 95238 76350
rect 95294 76294 95362 76350
rect 95418 76294 95488 76350
rect 95168 76226 95488 76294
rect 95168 76170 95238 76226
rect 95294 76170 95362 76226
rect 95418 76170 95488 76226
rect 95168 76102 95488 76170
rect 95168 76046 95238 76102
rect 95294 76046 95362 76102
rect 95418 76046 95488 76102
rect 95168 75978 95488 76046
rect 95168 75922 95238 75978
rect 95294 75922 95362 75978
rect 95418 75922 95488 75978
rect 95168 75888 95488 75922
rect 125888 76350 126208 76384
rect 125888 76294 125958 76350
rect 126014 76294 126082 76350
rect 126138 76294 126208 76350
rect 125888 76226 126208 76294
rect 125888 76170 125958 76226
rect 126014 76170 126082 76226
rect 126138 76170 126208 76226
rect 125888 76102 126208 76170
rect 125888 76046 125958 76102
rect 126014 76046 126082 76102
rect 126138 76046 126208 76102
rect 125888 75978 126208 76046
rect 125888 75922 125958 75978
rect 126014 75922 126082 75978
rect 126138 75922 126208 75978
rect 125888 75888 126208 75922
rect 156608 76350 156928 76384
rect 156608 76294 156678 76350
rect 156734 76294 156802 76350
rect 156858 76294 156928 76350
rect 156608 76226 156928 76294
rect 156608 76170 156678 76226
rect 156734 76170 156802 76226
rect 156858 76170 156928 76226
rect 156608 76102 156928 76170
rect 156608 76046 156678 76102
rect 156734 76046 156802 76102
rect 156858 76046 156928 76102
rect 156608 75978 156928 76046
rect 156608 75922 156678 75978
rect 156734 75922 156802 75978
rect 156858 75922 156928 75978
rect 156608 75888 156928 75922
rect 187328 76350 187648 76384
rect 187328 76294 187398 76350
rect 187454 76294 187522 76350
rect 187578 76294 187648 76350
rect 187328 76226 187648 76294
rect 187328 76170 187398 76226
rect 187454 76170 187522 76226
rect 187578 76170 187648 76226
rect 187328 76102 187648 76170
rect 187328 76046 187398 76102
rect 187454 76046 187522 76102
rect 187578 76046 187648 76102
rect 187328 75978 187648 76046
rect 187328 75922 187398 75978
rect 187454 75922 187522 75978
rect 187578 75922 187648 75978
rect 187328 75888 187648 75922
rect 218048 76350 218368 76384
rect 218048 76294 218118 76350
rect 218174 76294 218242 76350
rect 218298 76294 218368 76350
rect 218048 76226 218368 76294
rect 218048 76170 218118 76226
rect 218174 76170 218242 76226
rect 218298 76170 218368 76226
rect 218048 76102 218368 76170
rect 218048 76046 218118 76102
rect 218174 76046 218242 76102
rect 218298 76046 218368 76102
rect 218048 75978 218368 76046
rect 218048 75922 218118 75978
rect 218174 75922 218242 75978
rect 218298 75922 218368 75978
rect 218048 75888 218368 75922
rect 248768 76350 249088 76384
rect 248768 76294 248838 76350
rect 248894 76294 248962 76350
rect 249018 76294 249088 76350
rect 248768 76226 249088 76294
rect 248768 76170 248838 76226
rect 248894 76170 248962 76226
rect 249018 76170 249088 76226
rect 248768 76102 249088 76170
rect 248768 76046 248838 76102
rect 248894 76046 248962 76102
rect 249018 76046 249088 76102
rect 248768 75978 249088 76046
rect 248768 75922 248838 75978
rect 248894 75922 248962 75978
rect 249018 75922 249088 75978
rect 248768 75888 249088 75922
rect 279488 76350 279808 76384
rect 279488 76294 279558 76350
rect 279614 76294 279682 76350
rect 279738 76294 279808 76350
rect 279488 76226 279808 76294
rect 279488 76170 279558 76226
rect 279614 76170 279682 76226
rect 279738 76170 279808 76226
rect 279488 76102 279808 76170
rect 279488 76046 279558 76102
rect 279614 76046 279682 76102
rect 279738 76046 279808 76102
rect 279488 75978 279808 76046
rect 279488 75922 279558 75978
rect 279614 75922 279682 75978
rect 279738 75922 279808 75978
rect 279488 75888 279808 75922
rect 310208 76350 310528 76384
rect 310208 76294 310278 76350
rect 310334 76294 310402 76350
rect 310458 76294 310528 76350
rect 310208 76226 310528 76294
rect 310208 76170 310278 76226
rect 310334 76170 310402 76226
rect 310458 76170 310528 76226
rect 310208 76102 310528 76170
rect 310208 76046 310278 76102
rect 310334 76046 310402 76102
rect 310458 76046 310528 76102
rect 310208 75978 310528 76046
rect 310208 75922 310278 75978
rect 310334 75922 310402 75978
rect 310458 75922 310528 75978
rect 310208 75888 310528 75922
rect 340928 76350 341248 76384
rect 340928 76294 340998 76350
rect 341054 76294 341122 76350
rect 341178 76294 341248 76350
rect 340928 76226 341248 76294
rect 340928 76170 340998 76226
rect 341054 76170 341122 76226
rect 341178 76170 341248 76226
rect 340928 76102 341248 76170
rect 340928 76046 340998 76102
rect 341054 76046 341122 76102
rect 341178 76046 341248 76102
rect 340928 75978 341248 76046
rect 340928 75922 340998 75978
rect 341054 75922 341122 75978
rect 341178 75922 341248 75978
rect 340928 75888 341248 75922
rect 79808 64350 80128 64384
rect 79808 64294 79878 64350
rect 79934 64294 80002 64350
rect 80058 64294 80128 64350
rect 79808 64226 80128 64294
rect 79808 64170 79878 64226
rect 79934 64170 80002 64226
rect 80058 64170 80128 64226
rect 79808 64102 80128 64170
rect 79808 64046 79878 64102
rect 79934 64046 80002 64102
rect 80058 64046 80128 64102
rect 79808 63978 80128 64046
rect 79808 63922 79878 63978
rect 79934 63922 80002 63978
rect 80058 63922 80128 63978
rect 79808 63888 80128 63922
rect 110528 64350 110848 64384
rect 110528 64294 110598 64350
rect 110654 64294 110722 64350
rect 110778 64294 110848 64350
rect 110528 64226 110848 64294
rect 110528 64170 110598 64226
rect 110654 64170 110722 64226
rect 110778 64170 110848 64226
rect 110528 64102 110848 64170
rect 110528 64046 110598 64102
rect 110654 64046 110722 64102
rect 110778 64046 110848 64102
rect 110528 63978 110848 64046
rect 110528 63922 110598 63978
rect 110654 63922 110722 63978
rect 110778 63922 110848 63978
rect 110528 63888 110848 63922
rect 141248 64350 141568 64384
rect 141248 64294 141318 64350
rect 141374 64294 141442 64350
rect 141498 64294 141568 64350
rect 141248 64226 141568 64294
rect 141248 64170 141318 64226
rect 141374 64170 141442 64226
rect 141498 64170 141568 64226
rect 141248 64102 141568 64170
rect 141248 64046 141318 64102
rect 141374 64046 141442 64102
rect 141498 64046 141568 64102
rect 141248 63978 141568 64046
rect 141248 63922 141318 63978
rect 141374 63922 141442 63978
rect 141498 63922 141568 63978
rect 141248 63888 141568 63922
rect 171968 64350 172288 64384
rect 171968 64294 172038 64350
rect 172094 64294 172162 64350
rect 172218 64294 172288 64350
rect 171968 64226 172288 64294
rect 171968 64170 172038 64226
rect 172094 64170 172162 64226
rect 172218 64170 172288 64226
rect 171968 64102 172288 64170
rect 171968 64046 172038 64102
rect 172094 64046 172162 64102
rect 172218 64046 172288 64102
rect 171968 63978 172288 64046
rect 171968 63922 172038 63978
rect 172094 63922 172162 63978
rect 172218 63922 172288 63978
rect 171968 63888 172288 63922
rect 202688 64350 203008 64384
rect 202688 64294 202758 64350
rect 202814 64294 202882 64350
rect 202938 64294 203008 64350
rect 202688 64226 203008 64294
rect 202688 64170 202758 64226
rect 202814 64170 202882 64226
rect 202938 64170 203008 64226
rect 202688 64102 203008 64170
rect 202688 64046 202758 64102
rect 202814 64046 202882 64102
rect 202938 64046 203008 64102
rect 202688 63978 203008 64046
rect 202688 63922 202758 63978
rect 202814 63922 202882 63978
rect 202938 63922 203008 63978
rect 202688 63888 203008 63922
rect 233408 64350 233728 64384
rect 233408 64294 233478 64350
rect 233534 64294 233602 64350
rect 233658 64294 233728 64350
rect 233408 64226 233728 64294
rect 233408 64170 233478 64226
rect 233534 64170 233602 64226
rect 233658 64170 233728 64226
rect 233408 64102 233728 64170
rect 233408 64046 233478 64102
rect 233534 64046 233602 64102
rect 233658 64046 233728 64102
rect 233408 63978 233728 64046
rect 233408 63922 233478 63978
rect 233534 63922 233602 63978
rect 233658 63922 233728 63978
rect 233408 63888 233728 63922
rect 264128 64350 264448 64384
rect 264128 64294 264198 64350
rect 264254 64294 264322 64350
rect 264378 64294 264448 64350
rect 264128 64226 264448 64294
rect 264128 64170 264198 64226
rect 264254 64170 264322 64226
rect 264378 64170 264448 64226
rect 264128 64102 264448 64170
rect 264128 64046 264198 64102
rect 264254 64046 264322 64102
rect 264378 64046 264448 64102
rect 264128 63978 264448 64046
rect 264128 63922 264198 63978
rect 264254 63922 264322 63978
rect 264378 63922 264448 63978
rect 264128 63888 264448 63922
rect 294848 64350 295168 64384
rect 294848 64294 294918 64350
rect 294974 64294 295042 64350
rect 295098 64294 295168 64350
rect 294848 64226 295168 64294
rect 294848 64170 294918 64226
rect 294974 64170 295042 64226
rect 295098 64170 295168 64226
rect 294848 64102 295168 64170
rect 294848 64046 294918 64102
rect 294974 64046 295042 64102
rect 295098 64046 295168 64102
rect 294848 63978 295168 64046
rect 294848 63922 294918 63978
rect 294974 63922 295042 63978
rect 295098 63922 295168 63978
rect 294848 63888 295168 63922
rect 325568 64350 325888 64384
rect 325568 64294 325638 64350
rect 325694 64294 325762 64350
rect 325818 64294 325888 64350
rect 325568 64226 325888 64294
rect 325568 64170 325638 64226
rect 325694 64170 325762 64226
rect 325818 64170 325888 64226
rect 325568 64102 325888 64170
rect 325568 64046 325638 64102
rect 325694 64046 325762 64102
rect 325818 64046 325888 64102
rect 325568 63978 325888 64046
rect 325568 63922 325638 63978
rect 325694 63922 325762 63978
rect 325818 63922 325888 63978
rect 325568 63888 325888 63922
rect 348874 64350 349494 81922
rect 356288 82350 356608 82384
rect 356288 82294 356358 82350
rect 356414 82294 356482 82350
rect 356538 82294 356608 82350
rect 356288 82226 356608 82294
rect 356288 82170 356358 82226
rect 356414 82170 356482 82226
rect 356538 82170 356608 82226
rect 356288 82102 356608 82170
rect 356288 82046 356358 82102
rect 356414 82046 356482 82102
rect 356538 82046 356608 82102
rect 356288 81978 356608 82046
rect 356288 81922 356358 81978
rect 356414 81922 356482 81978
rect 356538 81922 356608 81978
rect 356288 81888 356608 81922
rect 363154 76350 363774 93922
rect 363154 76294 363250 76350
rect 363306 76294 363374 76350
rect 363430 76294 363498 76350
rect 363554 76294 363622 76350
rect 363678 76294 363774 76350
rect 363154 76226 363774 76294
rect 363154 76170 363250 76226
rect 363306 76170 363374 76226
rect 363430 76170 363498 76226
rect 363554 76170 363622 76226
rect 363678 76170 363774 76226
rect 363154 76102 363774 76170
rect 363154 76046 363250 76102
rect 363306 76046 363374 76102
rect 363430 76046 363498 76102
rect 363554 76046 363622 76102
rect 363678 76046 363774 76102
rect 363154 75978 363774 76046
rect 363154 75922 363250 75978
rect 363306 75922 363374 75978
rect 363430 75922 363498 75978
rect 363554 75922 363622 75978
rect 363678 75922 363774 75978
rect 348874 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 349494 64350
rect 348874 64226 349494 64294
rect 348874 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 349494 64226
rect 348874 64102 349494 64170
rect 348874 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 349494 64102
rect 348874 63978 349494 64046
rect 348874 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 349494 63978
rect 57154 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 57774 58350
rect 57154 58226 57774 58294
rect 57154 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 57774 58226
rect 57154 58102 57774 58170
rect 57154 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 57774 58102
rect 57154 57978 57774 58046
rect 57154 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 57774 57978
rect 57154 40350 57774 57922
rect 57154 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 57774 40350
rect 57154 40226 57774 40294
rect 57154 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 57774 40226
rect 57154 40102 57774 40170
rect 57154 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 57774 40102
rect 57154 39978 57774 40046
rect 57154 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 57774 39978
rect 57154 22350 57774 39922
rect 57154 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 57774 22350
rect 57154 22226 57774 22294
rect 57154 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 57774 22226
rect 57154 22102 57774 22170
rect 57154 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 57774 22102
rect 57154 21978 57774 22046
rect 57154 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 57774 21978
rect 57154 4350 57774 21922
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 46350 61494 59082
rect 60874 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 61494 46350
rect 60874 46226 61494 46294
rect 60874 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 61494 46226
rect 60874 46102 61494 46170
rect 60874 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 61494 46102
rect 60874 45978 61494 46046
rect 60874 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 61494 45978
rect 60874 28350 61494 45922
rect 60874 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 61494 28350
rect 60874 28226 61494 28294
rect 60874 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 61494 28226
rect 60874 28102 61494 28170
rect 60874 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 61494 28102
rect 60874 27978 61494 28046
rect 60874 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 61494 27978
rect 60874 10350 61494 27922
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 58350 75774 59082
rect 75154 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 75774 58350
rect 75154 58226 75774 58294
rect 75154 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 75774 58226
rect 75154 58102 75774 58170
rect 75154 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 75774 58102
rect 75154 57978 75774 58046
rect 75154 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 75774 57978
rect 75154 40350 75774 57922
rect 75154 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 75774 40350
rect 75154 40226 75774 40294
rect 75154 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 75774 40226
rect 75154 40102 75774 40170
rect 75154 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 75774 40102
rect 75154 39978 75774 40046
rect 75154 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 75774 39978
rect 75154 22350 75774 39922
rect 75154 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 75774 22350
rect 75154 22226 75774 22294
rect 75154 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 75774 22226
rect 75154 22102 75774 22170
rect 75154 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 75774 22102
rect 75154 21978 75774 22046
rect 75154 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 75774 21978
rect 75154 4350 75774 21922
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 46350 79494 59082
rect 78874 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 79494 46350
rect 78874 46226 79494 46294
rect 78874 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 79494 46226
rect 78874 46102 79494 46170
rect 78874 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 79494 46102
rect 78874 45978 79494 46046
rect 78874 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 79494 45978
rect 78874 28350 79494 45922
rect 78874 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 79494 28350
rect 78874 28226 79494 28294
rect 78874 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 79494 28226
rect 78874 28102 79494 28170
rect 78874 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 79494 28102
rect 78874 27978 79494 28046
rect 78874 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 79494 27978
rect 78874 10350 79494 27922
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 58350 93774 59082
rect 93154 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 93774 58350
rect 93154 58226 93774 58294
rect 93154 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 93774 58226
rect 93154 58102 93774 58170
rect 93154 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 93774 58102
rect 93154 57978 93774 58046
rect 93154 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 93774 57978
rect 93154 40350 93774 57922
rect 93154 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 93774 40350
rect 93154 40226 93774 40294
rect 93154 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 93774 40226
rect 93154 40102 93774 40170
rect 93154 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 93774 40102
rect 93154 39978 93774 40046
rect 93154 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 93774 39978
rect 93154 22350 93774 39922
rect 93154 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 93774 22350
rect 93154 22226 93774 22294
rect 93154 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 93774 22226
rect 93154 22102 93774 22170
rect 93154 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 93774 22102
rect 93154 21978 93774 22046
rect 93154 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 93774 21978
rect 93154 4350 93774 21922
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 46350 97494 59082
rect 96874 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 97494 46350
rect 96874 46226 97494 46294
rect 96874 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 97494 46226
rect 96874 46102 97494 46170
rect 96874 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 97494 46102
rect 96874 45978 97494 46046
rect 96874 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 97494 45978
rect 96874 28350 97494 45922
rect 96874 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 97494 28350
rect 96874 28226 97494 28294
rect 96874 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 97494 28226
rect 96874 28102 97494 28170
rect 96874 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 97494 28102
rect 96874 27978 97494 28046
rect 96874 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 97494 27978
rect 96874 10350 97494 27922
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 58350 111774 59082
rect 111154 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 111774 58350
rect 111154 58226 111774 58294
rect 111154 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 111774 58226
rect 111154 58102 111774 58170
rect 111154 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 111774 58102
rect 111154 57978 111774 58046
rect 111154 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 111774 57978
rect 111154 40350 111774 57922
rect 111154 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 111774 40350
rect 111154 40226 111774 40294
rect 111154 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 111774 40226
rect 111154 40102 111774 40170
rect 111154 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 111774 40102
rect 111154 39978 111774 40046
rect 111154 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 111774 39978
rect 111154 22350 111774 39922
rect 111154 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 111774 22350
rect 111154 22226 111774 22294
rect 111154 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 111774 22226
rect 111154 22102 111774 22170
rect 111154 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 111774 22102
rect 111154 21978 111774 22046
rect 111154 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 111774 21978
rect 111154 4350 111774 21922
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 46350 115494 59082
rect 114874 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 115494 46350
rect 114874 46226 115494 46294
rect 114874 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 115494 46226
rect 114874 46102 115494 46170
rect 114874 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 115494 46102
rect 114874 45978 115494 46046
rect 114874 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 115494 45978
rect 114874 28350 115494 45922
rect 114874 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 115494 28350
rect 114874 28226 115494 28294
rect 114874 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 115494 28226
rect 114874 28102 115494 28170
rect 114874 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 115494 28102
rect 114874 27978 115494 28046
rect 114874 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 115494 27978
rect 114874 10350 115494 27922
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 58350 129774 59082
rect 129154 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 129774 58350
rect 129154 58226 129774 58294
rect 129154 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 129774 58226
rect 129154 58102 129774 58170
rect 129154 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 129774 58102
rect 129154 57978 129774 58046
rect 129154 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 129774 57978
rect 129154 40350 129774 57922
rect 129154 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 129774 40350
rect 129154 40226 129774 40294
rect 129154 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 129774 40226
rect 129154 40102 129774 40170
rect 129154 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 129774 40102
rect 129154 39978 129774 40046
rect 129154 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 129774 39978
rect 129154 22350 129774 39922
rect 129154 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 129774 22350
rect 129154 22226 129774 22294
rect 129154 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 129774 22226
rect 129154 22102 129774 22170
rect 129154 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 129774 22102
rect 129154 21978 129774 22046
rect 129154 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 129774 21978
rect 129154 4350 129774 21922
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 46350 133494 59082
rect 132874 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 133494 46350
rect 132874 46226 133494 46294
rect 132874 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 133494 46226
rect 132874 46102 133494 46170
rect 132874 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 133494 46102
rect 132874 45978 133494 46046
rect 132874 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 133494 45978
rect 132874 28350 133494 45922
rect 132874 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 133494 28350
rect 132874 28226 133494 28294
rect 132874 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 133494 28226
rect 132874 28102 133494 28170
rect 132874 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 133494 28102
rect 132874 27978 133494 28046
rect 132874 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 133494 27978
rect 132874 10350 133494 27922
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 58350 147774 59082
rect 147154 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 147774 58350
rect 147154 58226 147774 58294
rect 147154 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 147774 58226
rect 147154 58102 147774 58170
rect 147154 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 147774 58102
rect 147154 57978 147774 58046
rect 147154 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 147774 57978
rect 147154 40350 147774 57922
rect 147154 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 147774 40350
rect 147154 40226 147774 40294
rect 147154 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 147774 40226
rect 147154 40102 147774 40170
rect 147154 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 147774 40102
rect 147154 39978 147774 40046
rect 147154 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 147774 39978
rect 147154 22350 147774 39922
rect 147154 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 147774 22350
rect 147154 22226 147774 22294
rect 147154 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 147774 22226
rect 147154 22102 147774 22170
rect 147154 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 147774 22102
rect 147154 21978 147774 22046
rect 147154 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 147774 21978
rect 147154 4350 147774 21922
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 46350 151494 59082
rect 150874 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 151494 46350
rect 150874 46226 151494 46294
rect 150874 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 151494 46226
rect 150874 46102 151494 46170
rect 150874 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 151494 46102
rect 150874 45978 151494 46046
rect 150874 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 151494 45978
rect 150874 28350 151494 45922
rect 150874 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 151494 28350
rect 150874 28226 151494 28294
rect 150874 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 151494 28226
rect 150874 28102 151494 28170
rect 150874 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 151494 28102
rect 150874 27978 151494 28046
rect 150874 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 151494 27978
rect 150874 10350 151494 27922
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 58350 165774 59082
rect 165154 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 165774 58350
rect 165154 58226 165774 58294
rect 165154 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 165774 58226
rect 165154 58102 165774 58170
rect 165154 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 165774 58102
rect 165154 57978 165774 58046
rect 165154 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 165774 57978
rect 165154 40350 165774 57922
rect 165154 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 165774 40350
rect 165154 40226 165774 40294
rect 165154 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 165774 40226
rect 165154 40102 165774 40170
rect 165154 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 165774 40102
rect 165154 39978 165774 40046
rect 165154 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 165774 39978
rect 165154 22350 165774 39922
rect 165154 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 165774 22350
rect 165154 22226 165774 22294
rect 165154 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 165774 22226
rect 165154 22102 165774 22170
rect 165154 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 165774 22102
rect 165154 21978 165774 22046
rect 165154 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 165774 21978
rect 165154 4350 165774 21922
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 46350 169494 59082
rect 168874 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 169494 46350
rect 168874 46226 169494 46294
rect 168874 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 169494 46226
rect 168874 46102 169494 46170
rect 168874 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 169494 46102
rect 168874 45978 169494 46046
rect 168874 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 169494 45978
rect 168874 28350 169494 45922
rect 168874 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 169494 28350
rect 168874 28226 169494 28294
rect 168874 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 169494 28226
rect 168874 28102 169494 28170
rect 168874 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 169494 28102
rect 168874 27978 169494 28046
rect 168874 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 169494 27978
rect 168874 10350 169494 27922
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 58350 183774 59082
rect 183154 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 183774 58350
rect 183154 58226 183774 58294
rect 183154 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 183774 58226
rect 183154 58102 183774 58170
rect 183154 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 183774 58102
rect 183154 57978 183774 58046
rect 183154 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 183774 57978
rect 183154 40350 183774 57922
rect 183154 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 183774 40350
rect 183154 40226 183774 40294
rect 183154 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 183774 40226
rect 183154 40102 183774 40170
rect 183154 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 183774 40102
rect 183154 39978 183774 40046
rect 183154 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 183774 39978
rect 183154 22350 183774 39922
rect 183154 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 183774 22350
rect 183154 22226 183774 22294
rect 183154 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 183774 22226
rect 183154 22102 183774 22170
rect 183154 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 183774 22102
rect 183154 21978 183774 22046
rect 183154 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 183774 21978
rect 183154 4350 183774 21922
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 46350 187494 59082
rect 186874 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 187494 46350
rect 186874 46226 187494 46294
rect 186874 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 187494 46226
rect 186874 46102 187494 46170
rect 186874 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 187494 46102
rect 186874 45978 187494 46046
rect 186874 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 187494 45978
rect 186874 28350 187494 45922
rect 186874 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 187494 28350
rect 186874 28226 187494 28294
rect 186874 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 187494 28226
rect 186874 28102 187494 28170
rect 186874 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 187494 28102
rect 186874 27978 187494 28046
rect 186874 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 187494 27978
rect 186874 10350 187494 27922
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 58350 201774 59082
rect 201154 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 201774 58350
rect 201154 58226 201774 58294
rect 201154 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 201774 58226
rect 201154 58102 201774 58170
rect 201154 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 201774 58102
rect 201154 57978 201774 58046
rect 201154 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 201774 57978
rect 201154 40350 201774 57922
rect 201154 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 201774 40350
rect 201154 40226 201774 40294
rect 201154 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 201774 40226
rect 201154 40102 201774 40170
rect 201154 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 201774 40102
rect 201154 39978 201774 40046
rect 201154 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 201774 39978
rect 201154 22350 201774 39922
rect 201154 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 201774 22350
rect 201154 22226 201774 22294
rect 201154 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 201774 22226
rect 201154 22102 201774 22170
rect 201154 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 201774 22102
rect 201154 21978 201774 22046
rect 201154 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 201774 21978
rect 201154 4350 201774 21922
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 46350 205494 59082
rect 204874 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 205494 46350
rect 204874 46226 205494 46294
rect 204874 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 205494 46226
rect 204874 46102 205494 46170
rect 204874 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 205494 46102
rect 204874 45978 205494 46046
rect 204874 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 205494 45978
rect 204874 28350 205494 45922
rect 204874 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 205494 28350
rect 204874 28226 205494 28294
rect 204874 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 205494 28226
rect 204874 28102 205494 28170
rect 204874 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 205494 28102
rect 204874 27978 205494 28046
rect 204874 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 205494 27978
rect 204874 10350 205494 27922
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 58350 219774 59082
rect 219154 58294 219250 58350
rect 219306 58294 219374 58350
rect 219430 58294 219498 58350
rect 219554 58294 219622 58350
rect 219678 58294 219774 58350
rect 219154 58226 219774 58294
rect 219154 58170 219250 58226
rect 219306 58170 219374 58226
rect 219430 58170 219498 58226
rect 219554 58170 219622 58226
rect 219678 58170 219774 58226
rect 219154 58102 219774 58170
rect 219154 58046 219250 58102
rect 219306 58046 219374 58102
rect 219430 58046 219498 58102
rect 219554 58046 219622 58102
rect 219678 58046 219774 58102
rect 219154 57978 219774 58046
rect 219154 57922 219250 57978
rect 219306 57922 219374 57978
rect 219430 57922 219498 57978
rect 219554 57922 219622 57978
rect 219678 57922 219774 57978
rect 219154 40350 219774 57922
rect 219154 40294 219250 40350
rect 219306 40294 219374 40350
rect 219430 40294 219498 40350
rect 219554 40294 219622 40350
rect 219678 40294 219774 40350
rect 219154 40226 219774 40294
rect 219154 40170 219250 40226
rect 219306 40170 219374 40226
rect 219430 40170 219498 40226
rect 219554 40170 219622 40226
rect 219678 40170 219774 40226
rect 219154 40102 219774 40170
rect 219154 40046 219250 40102
rect 219306 40046 219374 40102
rect 219430 40046 219498 40102
rect 219554 40046 219622 40102
rect 219678 40046 219774 40102
rect 219154 39978 219774 40046
rect 219154 39922 219250 39978
rect 219306 39922 219374 39978
rect 219430 39922 219498 39978
rect 219554 39922 219622 39978
rect 219678 39922 219774 39978
rect 219154 22350 219774 39922
rect 219154 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 219774 22350
rect 219154 22226 219774 22294
rect 219154 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 219774 22226
rect 219154 22102 219774 22170
rect 219154 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 219774 22102
rect 219154 21978 219774 22046
rect 219154 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 219774 21978
rect 219154 4350 219774 21922
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 222874 46350 223494 59082
rect 222874 46294 222970 46350
rect 223026 46294 223094 46350
rect 223150 46294 223218 46350
rect 223274 46294 223342 46350
rect 223398 46294 223494 46350
rect 222874 46226 223494 46294
rect 222874 46170 222970 46226
rect 223026 46170 223094 46226
rect 223150 46170 223218 46226
rect 223274 46170 223342 46226
rect 223398 46170 223494 46226
rect 222874 46102 223494 46170
rect 222874 46046 222970 46102
rect 223026 46046 223094 46102
rect 223150 46046 223218 46102
rect 223274 46046 223342 46102
rect 223398 46046 223494 46102
rect 222874 45978 223494 46046
rect 222874 45922 222970 45978
rect 223026 45922 223094 45978
rect 223150 45922 223218 45978
rect 223274 45922 223342 45978
rect 223398 45922 223494 45978
rect 222874 28350 223494 45922
rect 222874 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 223494 28350
rect 222874 28226 223494 28294
rect 222874 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 223494 28226
rect 222874 28102 223494 28170
rect 222874 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 223494 28102
rect 222874 27978 223494 28046
rect 222874 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 223494 27978
rect 222874 10350 223494 27922
rect 222874 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 223494 10350
rect 222874 10226 223494 10294
rect 222874 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 223494 10226
rect 222874 10102 223494 10170
rect 222874 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 223494 10102
rect 222874 9978 223494 10046
rect 222874 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 223494 9978
rect 222874 -1120 223494 9922
rect 222874 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 223494 -1120
rect 222874 -1244 223494 -1176
rect 222874 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 223494 -1244
rect 222874 -1368 223494 -1300
rect 222874 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 223494 -1368
rect 222874 -1492 223494 -1424
rect 222874 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 223494 -1492
rect 222874 -1644 223494 -1548
rect 237154 58350 237774 59082
rect 237154 58294 237250 58350
rect 237306 58294 237374 58350
rect 237430 58294 237498 58350
rect 237554 58294 237622 58350
rect 237678 58294 237774 58350
rect 237154 58226 237774 58294
rect 237154 58170 237250 58226
rect 237306 58170 237374 58226
rect 237430 58170 237498 58226
rect 237554 58170 237622 58226
rect 237678 58170 237774 58226
rect 237154 58102 237774 58170
rect 237154 58046 237250 58102
rect 237306 58046 237374 58102
rect 237430 58046 237498 58102
rect 237554 58046 237622 58102
rect 237678 58046 237774 58102
rect 237154 57978 237774 58046
rect 237154 57922 237250 57978
rect 237306 57922 237374 57978
rect 237430 57922 237498 57978
rect 237554 57922 237622 57978
rect 237678 57922 237774 57978
rect 237154 40350 237774 57922
rect 237154 40294 237250 40350
rect 237306 40294 237374 40350
rect 237430 40294 237498 40350
rect 237554 40294 237622 40350
rect 237678 40294 237774 40350
rect 237154 40226 237774 40294
rect 237154 40170 237250 40226
rect 237306 40170 237374 40226
rect 237430 40170 237498 40226
rect 237554 40170 237622 40226
rect 237678 40170 237774 40226
rect 237154 40102 237774 40170
rect 237154 40046 237250 40102
rect 237306 40046 237374 40102
rect 237430 40046 237498 40102
rect 237554 40046 237622 40102
rect 237678 40046 237774 40102
rect 237154 39978 237774 40046
rect 237154 39922 237250 39978
rect 237306 39922 237374 39978
rect 237430 39922 237498 39978
rect 237554 39922 237622 39978
rect 237678 39922 237774 39978
rect 237154 22350 237774 39922
rect 237154 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 237774 22350
rect 237154 22226 237774 22294
rect 237154 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 237774 22226
rect 237154 22102 237774 22170
rect 237154 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 237774 22102
rect 237154 21978 237774 22046
rect 237154 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 237774 21978
rect 237154 4350 237774 21922
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 240874 46350 241494 59082
rect 240874 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 241494 46350
rect 240874 46226 241494 46294
rect 240874 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 241494 46226
rect 240874 46102 241494 46170
rect 240874 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 241494 46102
rect 240874 45978 241494 46046
rect 240874 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 241494 45978
rect 240874 28350 241494 45922
rect 240874 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 241494 28350
rect 240874 28226 241494 28294
rect 240874 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 241494 28226
rect 240874 28102 241494 28170
rect 240874 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 241494 28102
rect 240874 27978 241494 28046
rect 240874 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 241494 27978
rect 240874 10350 241494 27922
rect 240874 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 241494 10350
rect 240874 10226 241494 10294
rect 240874 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 241494 10226
rect 240874 10102 241494 10170
rect 240874 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 241494 10102
rect 240874 9978 241494 10046
rect 240874 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 241494 9978
rect 240874 -1120 241494 9922
rect 240874 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 241494 -1120
rect 240874 -1244 241494 -1176
rect 240874 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 241494 -1244
rect 240874 -1368 241494 -1300
rect 240874 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 241494 -1368
rect 240874 -1492 241494 -1424
rect 240874 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 241494 -1492
rect 240874 -1644 241494 -1548
rect 255154 58350 255774 59082
rect 255154 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 255774 58350
rect 255154 58226 255774 58294
rect 255154 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 255774 58226
rect 255154 58102 255774 58170
rect 255154 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 255774 58102
rect 255154 57978 255774 58046
rect 255154 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 255774 57978
rect 255154 40350 255774 57922
rect 255154 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 255774 40350
rect 255154 40226 255774 40294
rect 255154 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 255774 40226
rect 255154 40102 255774 40170
rect 255154 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 255774 40102
rect 255154 39978 255774 40046
rect 255154 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 255774 39978
rect 255154 22350 255774 39922
rect 255154 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 255774 22350
rect 255154 22226 255774 22294
rect 255154 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 255774 22226
rect 255154 22102 255774 22170
rect 255154 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 255774 22102
rect 255154 21978 255774 22046
rect 255154 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 255774 21978
rect 255154 4350 255774 21922
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 258874 46350 259494 59082
rect 258874 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 259494 46350
rect 258874 46226 259494 46294
rect 258874 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 259494 46226
rect 258874 46102 259494 46170
rect 258874 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 259494 46102
rect 258874 45978 259494 46046
rect 258874 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 259494 45978
rect 258874 28350 259494 45922
rect 258874 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 259494 28350
rect 258874 28226 259494 28294
rect 258874 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 259494 28226
rect 258874 28102 259494 28170
rect 258874 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 259494 28102
rect 258874 27978 259494 28046
rect 258874 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 259494 27978
rect 258874 10350 259494 27922
rect 258874 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 259494 10350
rect 258874 10226 259494 10294
rect 258874 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 259494 10226
rect 258874 10102 259494 10170
rect 258874 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 259494 10102
rect 258874 9978 259494 10046
rect 258874 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 259494 9978
rect 258874 -1120 259494 9922
rect 258874 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 259494 -1120
rect 258874 -1244 259494 -1176
rect 258874 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 259494 -1244
rect 258874 -1368 259494 -1300
rect 258874 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 259494 -1368
rect 258874 -1492 259494 -1424
rect 258874 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 259494 -1492
rect 258874 -1644 259494 -1548
rect 273154 58350 273774 59082
rect 273154 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 273774 58350
rect 273154 58226 273774 58294
rect 273154 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 273774 58226
rect 273154 58102 273774 58170
rect 273154 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 273774 58102
rect 273154 57978 273774 58046
rect 273154 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 273774 57978
rect 273154 40350 273774 57922
rect 273154 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 273774 40350
rect 273154 40226 273774 40294
rect 273154 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 273774 40226
rect 273154 40102 273774 40170
rect 273154 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 273774 40102
rect 273154 39978 273774 40046
rect 273154 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 273774 39978
rect 273154 22350 273774 39922
rect 273154 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 273774 22350
rect 273154 22226 273774 22294
rect 273154 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 273774 22226
rect 273154 22102 273774 22170
rect 273154 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 273774 22102
rect 273154 21978 273774 22046
rect 273154 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 273774 21978
rect 273154 4350 273774 21922
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 276874 46350 277494 59082
rect 276874 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 277494 46350
rect 276874 46226 277494 46294
rect 276874 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 277494 46226
rect 276874 46102 277494 46170
rect 276874 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 277494 46102
rect 276874 45978 277494 46046
rect 276874 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 277494 45978
rect 276874 28350 277494 45922
rect 276874 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 277494 28350
rect 276874 28226 277494 28294
rect 276874 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 277494 28226
rect 276874 28102 277494 28170
rect 276874 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 277494 28102
rect 276874 27978 277494 28046
rect 276874 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 277494 27978
rect 276874 10350 277494 27922
rect 276874 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 277494 10350
rect 276874 10226 277494 10294
rect 276874 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 277494 10226
rect 276874 10102 277494 10170
rect 276874 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 277494 10102
rect 276874 9978 277494 10046
rect 276874 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 277494 9978
rect 276874 -1120 277494 9922
rect 276874 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 277494 -1120
rect 276874 -1244 277494 -1176
rect 276874 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 277494 -1244
rect 276874 -1368 277494 -1300
rect 276874 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 277494 -1368
rect 276874 -1492 277494 -1424
rect 276874 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 277494 -1492
rect 276874 -1644 277494 -1548
rect 291154 58350 291774 59082
rect 291154 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 291774 58350
rect 291154 58226 291774 58294
rect 291154 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 291774 58226
rect 291154 58102 291774 58170
rect 291154 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 291774 58102
rect 291154 57978 291774 58046
rect 291154 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 291774 57978
rect 291154 40350 291774 57922
rect 291154 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 291774 40350
rect 291154 40226 291774 40294
rect 291154 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 291774 40226
rect 291154 40102 291774 40170
rect 291154 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 291774 40102
rect 291154 39978 291774 40046
rect 291154 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 291774 39978
rect 291154 22350 291774 39922
rect 291154 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 291774 22350
rect 291154 22226 291774 22294
rect 291154 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 291774 22226
rect 291154 22102 291774 22170
rect 291154 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 291774 22102
rect 291154 21978 291774 22046
rect 291154 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 291774 21978
rect 291154 4350 291774 21922
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 294874 46350 295494 59082
rect 294874 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 295494 46350
rect 294874 46226 295494 46294
rect 294874 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 295494 46226
rect 294874 46102 295494 46170
rect 294874 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 295494 46102
rect 294874 45978 295494 46046
rect 294874 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 295494 45978
rect 294874 28350 295494 45922
rect 294874 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 295494 28350
rect 294874 28226 295494 28294
rect 294874 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 295494 28226
rect 294874 28102 295494 28170
rect 294874 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 295494 28102
rect 294874 27978 295494 28046
rect 294874 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 295494 27978
rect 294874 10350 295494 27922
rect 294874 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 295494 10350
rect 294874 10226 295494 10294
rect 294874 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 295494 10226
rect 294874 10102 295494 10170
rect 294874 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 295494 10102
rect 294874 9978 295494 10046
rect 294874 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 295494 9978
rect 294874 -1120 295494 9922
rect 294874 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 295494 -1120
rect 294874 -1244 295494 -1176
rect 294874 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 295494 -1244
rect 294874 -1368 295494 -1300
rect 294874 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 295494 -1368
rect 294874 -1492 295494 -1424
rect 294874 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 295494 -1492
rect 294874 -1644 295494 -1548
rect 309154 58350 309774 59082
rect 309154 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 309774 58350
rect 309154 58226 309774 58294
rect 309154 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 309774 58226
rect 309154 58102 309774 58170
rect 309154 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 309774 58102
rect 309154 57978 309774 58046
rect 309154 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 309774 57978
rect 309154 40350 309774 57922
rect 309154 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 309774 40350
rect 309154 40226 309774 40294
rect 309154 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 309774 40226
rect 309154 40102 309774 40170
rect 309154 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 309774 40102
rect 309154 39978 309774 40046
rect 309154 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 309774 39978
rect 309154 22350 309774 39922
rect 309154 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 309774 22350
rect 309154 22226 309774 22294
rect 309154 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 309774 22226
rect 309154 22102 309774 22170
rect 309154 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 309774 22102
rect 309154 21978 309774 22046
rect 309154 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 309774 21978
rect 309154 4350 309774 21922
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 312874 46350 313494 59082
rect 312874 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 313494 46350
rect 312874 46226 313494 46294
rect 312874 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 313494 46226
rect 312874 46102 313494 46170
rect 312874 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 313494 46102
rect 312874 45978 313494 46046
rect 312874 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 313494 45978
rect 312874 28350 313494 45922
rect 312874 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 313494 28350
rect 312874 28226 313494 28294
rect 312874 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 313494 28226
rect 312874 28102 313494 28170
rect 312874 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 313494 28102
rect 312874 27978 313494 28046
rect 312874 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 313494 27978
rect 312874 10350 313494 27922
rect 312874 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 313494 10350
rect 312874 10226 313494 10294
rect 312874 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 313494 10226
rect 312874 10102 313494 10170
rect 312874 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 313494 10102
rect 312874 9978 313494 10046
rect 312874 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 313494 9978
rect 312874 -1120 313494 9922
rect 312874 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 313494 -1120
rect 312874 -1244 313494 -1176
rect 312874 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 313494 -1244
rect 312874 -1368 313494 -1300
rect 312874 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 313494 -1368
rect 312874 -1492 313494 -1424
rect 312874 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 313494 -1492
rect 312874 -1644 313494 -1548
rect 327154 58350 327774 59082
rect 327154 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 327774 58350
rect 327154 58226 327774 58294
rect 327154 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 327774 58226
rect 327154 58102 327774 58170
rect 327154 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 327774 58102
rect 327154 57978 327774 58046
rect 327154 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 327774 57978
rect 327154 40350 327774 57922
rect 327154 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 327774 40350
rect 327154 40226 327774 40294
rect 327154 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 327774 40226
rect 327154 40102 327774 40170
rect 327154 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 327774 40102
rect 327154 39978 327774 40046
rect 327154 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 327774 39978
rect 327154 22350 327774 39922
rect 327154 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 327774 22350
rect 327154 22226 327774 22294
rect 327154 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 327774 22226
rect 327154 22102 327774 22170
rect 327154 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 327774 22102
rect 327154 21978 327774 22046
rect 327154 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 327774 21978
rect 327154 4350 327774 21922
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 330874 46350 331494 59082
rect 330874 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 331494 46350
rect 330874 46226 331494 46294
rect 330874 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 331494 46226
rect 330874 46102 331494 46170
rect 330874 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 331494 46102
rect 330874 45978 331494 46046
rect 330874 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 331494 45978
rect 330874 28350 331494 45922
rect 330874 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 331494 28350
rect 330874 28226 331494 28294
rect 330874 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 331494 28226
rect 330874 28102 331494 28170
rect 330874 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 331494 28102
rect 330874 27978 331494 28046
rect 330874 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 331494 27978
rect 330874 10350 331494 27922
rect 330874 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 331494 10350
rect 330874 10226 331494 10294
rect 330874 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 331494 10226
rect 330874 10102 331494 10170
rect 330874 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 331494 10102
rect 330874 9978 331494 10046
rect 330874 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 331494 9978
rect 330874 -1120 331494 9922
rect 330874 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 331494 -1120
rect 330874 -1244 331494 -1176
rect 330874 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 331494 -1244
rect 330874 -1368 331494 -1300
rect 330874 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 331494 -1368
rect 330874 -1492 331494 -1424
rect 330874 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 331494 -1492
rect 330874 -1644 331494 -1548
rect 345154 58350 345774 59082
rect 345154 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 345774 58350
rect 345154 58226 345774 58294
rect 345154 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 345774 58226
rect 345154 58102 345774 58170
rect 345154 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 345774 58102
rect 345154 57978 345774 58046
rect 345154 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 345774 57978
rect 345154 40350 345774 57922
rect 345154 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 345774 40350
rect 345154 40226 345774 40294
rect 345154 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 345774 40226
rect 345154 40102 345774 40170
rect 345154 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 345774 40102
rect 345154 39978 345774 40046
rect 345154 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 345774 39978
rect 345154 22350 345774 39922
rect 345154 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 345774 22350
rect 345154 22226 345774 22294
rect 345154 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 345774 22226
rect 345154 22102 345774 22170
rect 345154 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 345774 22102
rect 345154 21978 345774 22046
rect 345154 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 345774 21978
rect 345154 4350 345774 21922
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 348874 46350 349494 63922
rect 356288 64350 356608 64384
rect 356288 64294 356358 64350
rect 356414 64294 356482 64350
rect 356538 64294 356608 64350
rect 356288 64226 356608 64294
rect 356288 64170 356358 64226
rect 356414 64170 356482 64226
rect 356538 64170 356608 64226
rect 356288 64102 356608 64170
rect 356288 64046 356358 64102
rect 356414 64046 356482 64102
rect 356538 64046 356608 64102
rect 356288 63978 356608 64046
rect 356288 63922 356358 63978
rect 356414 63922 356482 63978
rect 356538 63922 356608 63978
rect 356288 63888 356608 63922
rect 348874 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 349494 46350
rect 348874 46226 349494 46294
rect 348874 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 349494 46226
rect 348874 46102 349494 46170
rect 348874 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 349494 46102
rect 348874 45978 349494 46046
rect 348874 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 349494 45978
rect 348874 28350 349494 45922
rect 348874 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 349494 28350
rect 348874 28226 349494 28294
rect 348874 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 349494 28226
rect 348874 28102 349494 28170
rect 348874 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 349494 28102
rect 348874 27978 349494 28046
rect 348874 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 349494 27978
rect 348874 10350 349494 27922
rect 348874 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 349494 10350
rect 348874 10226 349494 10294
rect 348874 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 349494 10226
rect 348874 10102 349494 10170
rect 348874 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 349494 10102
rect 348874 9978 349494 10046
rect 348874 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 349494 9978
rect 348874 -1120 349494 9922
rect 348874 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 349494 -1120
rect 348874 -1244 349494 -1176
rect 348874 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 349494 -1244
rect 348874 -1368 349494 -1300
rect 348874 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 349494 -1368
rect 348874 -1492 349494 -1424
rect 348874 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 349494 -1492
rect 348874 -1644 349494 -1548
rect 363154 58350 363774 75922
rect 363154 58294 363250 58350
rect 363306 58294 363374 58350
rect 363430 58294 363498 58350
rect 363554 58294 363622 58350
rect 363678 58294 363774 58350
rect 363154 58226 363774 58294
rect 363154 58170 363250 58226
rect 363306 58170 363374 58226
rect 363430 58170 363498 58226
rect 363554 58170 363622 58226
rect 363678 58170 363774 58226
rect 363154 58102 363774 58170
rect 363154 58046 363250 58102
rect 363306 58046 363374 58102
rect 363430 58046 363498 58102
rect 363554 58046 363622 58102
rect 363678 58046 363774 58102
rect 363154 57978 363774 58046
rect 363154 57922 363250 57978
rect 363306 57922 363374 57978
rect 363430 57922 363498 57978
rect 363554 57922 363622 57978
rect 363678 57922 363774 57978
rect 363154 40350 363774 57922
rect 363154 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 363774 40350
rect 363154 40226 363774 40294
rect 363154 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 363774 40226
rect 363154 40102 363774 40170
rect 363154 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 363774 40102
rect 363154 39978 363774 40046
rect 363154 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 363774 39978
rect 363154 22350 363774 39922
rect 363154 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 363774 22350
rect 363154 22226 363774 22294
rect 363154 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 363774 22226
rect 363154 22102 363774 22170
rect 363154 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 363774 22102
rect 363154 21978 363774 22046
rect 363154 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 363774 21978
rect 363154 4350 363774 21922
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 514350 367494 531922
rect 366874 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 367494 514350
rect 366874 514226 367494 514294
rect 366874 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 367494 514226
rect 366874 514102 367494 514170
rect 366874 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 367494 514102
rect 366874 513978 367494 514046
rect 366874 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 367494 513978
rect 366874 496350 367494 513922
rect 366874 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 367494 496350
rect 366874 496226 367494 496294
rect 366874 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 367494 496226
rect 366874 496102 367494 496170
rect 366874 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 367494 496102
rect 366874 495978 367494 496046
rect 366874 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 367494 495978
rect 366874 478350 367494 495922
rect 366874 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 367494 478350
rect 366874 478226 367494 478294
rect 366874 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 367494 478226
rect 366874 478102 367494 478170
rect 366874 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 367494 478102
rect 366874 477978 367494 478046
rect 366874 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 367494 477978
rect 366874 460350 367494 477922
rect 366874 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 367494 460350
rect 366874 460226 367494 460294
rect 366874 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 367494 460226
rect 366874 460102 367494 460170
rect 366874 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 367494 460102
rect 366874 459978 367494 460046
rect 366874 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 367494 459978
rect 366874 442350 367494 459922
rect 366874 442294 366970 442350
rect 367026 442294 367094 442350
rect 367150 442294 367218 442350
rect 367274 442294 367342 442350
rect 367398 442294 367494 442350
rect 366874 442226 367494 442294
rect 366874 442170 366970 442226
rect 367026 442170 367094 442226
rect 367150 442170 367218 442226
rect 367274 442170 367342 442226
rect 367398 442170 367494 442226
rect 366874 442102 367494 442170
rect 366874 442046 366970 442102
rect 367026 442046 367094 442102
rect 367150 442046 367218 442102
rect 367274 442046 367342 442102
rect 367398 442046 367494 442102
rect 366874 441978 367494 442046
rect 366874 441922 366970 441978
rect 367026 441922 367094 441978
rect 367150 441922 367218 441978
rect 367274 441922 367342 441978
rect 367398 441922 367494 441978
rect 366874 424350 367494 441922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 526350 381774 543922
rect 381154 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 381774 526350
rect 381154 526226 381774 526294
rect 381154 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 381774 526226
rect 381154 526102 381774 526170
rect 381154 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 381774 526102
rect 381154 525978 381774 526046
rect 381154 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 381774 525978
rect 381154 508350 381774 525922
rect 381154 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 381774 508350
rect 381154 508226 381774 508294
rect 381154 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 381774 508226
rect 381154 508102 381774 508170
rect 381154 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 381774 508102
rect 381154 507978 381774 508046
rect 381154 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 381774 507978
rect 381154 490350 381774 507922
rect 381154 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 381774 490350
rect 381154 490226 381774 490294
rect 381154 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 381774 490226
rect 381154 490102 381774 490170
rect 381154 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 381774 490102
rect 381154 489978 381774 490046
rect 381154 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 381774 489978
rect 381154 472350 381774 489922
rect 381154 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 381774 472350
rect 381154 472226 381774 472294
rect 381154 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 381774 472226
rect 381154 472102 381774 472170
rect 381154 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 381774 472102
rect 381154 471978 381774 472046
rect 381154 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 381774 471978
rect 381154 454350 381774 471922
rect 381154 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 381774 454350
rect 381154 454226 381774 454294
rect 381154 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 381774 454226
rect 381154 454102 381774 454170
rect 381154 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 381774 454102
rect 381154 453978 381774 454046
rect 381154 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 381774 453978
rect 371648 436317 371968 436380
rect 371648 436261 371718 436317
rect 371774 436261 371842 436317
rect 371898 436261 371968 436317
rect 371648 436193 371968 436261
rect 371648 436137 371718 436193
rect 371774 436137 371842 436193
rect 371898 436137 371968 436193
rect 371648 436069 371968 436137
rect 371648 436013 371718 436069
rect 371774 436013 371842 436069
rect 371898 436013 371968 436069
rect 371648 435945 371968 436013
rect 371648 435889 371718 435945
rect 371774 435889 371842 435945
rect 371898 435889 371968 435945
rect 371648 435826 371968 435889
rect 381154 436350 381774 453922
rect 381154 436294 381250 436350
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 381774 436350
rect 381154 436226 381774 436294
rect 381154 436170 381250 436226
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 381774 436226
rect 381154 436102 381774 436170
rect 381154 436046 381250 436102
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 381774 436102
rect 381154 435978 381774 436046
rect 381154 435922 381250 435978
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 381774 435978
rect 366874 424294 366970 424350
rect 367026 424294 367094 424350
rect 367150 424294 367218 424350
rect 367274 424294 367342 424350
rect 367398 424294 367494 424350
rect 366874 424226 367494 424294
rect 366874 424170 366970 424226
rect 367026 424170 367094 424226
rect 367150 424170 367218 424226
rect 367274 424170 367342 424226
rect 367398 424170 367494 424226
rect 366874 424102 367494 424170
rect 366874 424046 366970 424102
rect 367026 424046 367094 424102
rect 367150 424046 367218 424102
rect 367274 424046 367342 424102
rect 367398 424046 367494 424102
rect 366874 423978 367494 424046
rect 366874 423922 366970 423978
rect 367026 423922 367094 423978
rect 367150 423922 367218 423978
rect 367274 423922 367342 423978
rect 367398 423922 367494 423978
rect 366874 406350 367494 423922
rect 371648 418350 371968 418384
rect 371648 418294 371718 418350
rect 371774 418294 371842 418350
rect 371898 418294 371968 418350
rect 371648 418226 371968 418294
rect 371648 418170 371718 418226
rect 371774 418170 371842 418226
rect 371898 418170 371968 418226
rect 371648 418102 371968 418170
rect 371648 418046 371718 418102
rect 371774 418046 371842 418102
rect 371898 418046 371968 418102
rect 371648 417978 371968 418046
rect 371648 417922 371718 417978
rect 371774 417922 371842 417978
rect 371898 417922 371968 417978
rect 371648 417888 371968 417922
rect 381154 418350 381774 435922
rect 381154 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 381774 418350
rect 381154 418226 381774 418294
rect 381154 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 381774 418226
rect 381154 418102 381774 418170
rect 381154 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 381774 418102
rect 381154 417978 381774 418046
rect 381154 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 381774 417978
rect 366874 406294 366970 406350
rect 367026 406294 367094 406350
rect 367150 406294 367218 406350
rect 367274 406294 367342 406350
rect 367398 406294 367494 406350
rect 366874 406226 367494 406294
rect 366874 406170 366970 406226
rect 367026 406170 367094 406226
rect 367150 406170 367218 406226
rect 367274 406170 367342 406226
rect 367398 406170 367494 406226
rect 366874 406102 367494 406170
rect 366874 406046 366970 406102
rect 367026 406046 367094 406102
rect 367150 406046 367218 406102
rect 367274 406046 367342 406102
rect 367398 406046 367494 406102
rect 366874 405978 367494 406046
rect 366874 405922 366970 405978
rect 367026 405922 367094 405978
rect 367150 405922 367218 405978
rect 367274 405922 367342 405978
rect 367398 405922 367494 405978
rect 366874 388350 367494 405922
rect 371648 400350 371968 400384
rect 371648 400294 371718 400350
rect 371774 400294 371842 400350
rect 371898 400294 371968 400350
rect 371648 400226 371968 400294
rect 371648 400170 371718 400226
rect 371774 400170 371842 400226
rect 371898 400170 371968 400226
rect 371648 400102 371968 400170
rect 371648 400046 371718 400102
rect 371774 400046 371842 400102
rect 371898 400046 371968 400102
rect 371648 399978 371968 400046
rect 371648 399922 371718 399978
rect 371774 399922 371842 399978
rect 371898 399922 371968 399978
rect 371648 399888 371968 399922
rect 381154 400350 381774 417922
rect 381154 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 381774 400350
rect 381154 400226 381774 400294
rect 381154 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 381774 400226
rect 381154 400102 381774 400170
rect 381154 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 381774 400102
rect 381154 399978 381774 400046
rect 381154 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 381774 399978
rect 366874 388294 366970 388350
rect 367026 388294 367094 388350
rect 367150 388294 367218 388350
rect 367274 388294 367342 388350
rect 367398 388294 367494 388350
rect 366874 388226 367494 388294
rect 366874 388170 366970 388226
rect 367026 388170 367094 388226
rect 367150 388170 367218 388226
rect 367274 388170 367342 388226
rect 367398 388170 367494 388226
rect 366874 388102 367494 388170
rect 366874 388046 366970 388102
rect 367026 388046 367094 388102
rect 367150 388046 367218 388102
rect 367274 388046 367342 388102
rect 367398 388046 367494 388102
rect 366874 387978 367494 388046
rect 366874 387922 366970 387978
rect 367026 387922 367094 387978
rect 367150 387922 367218 387978
rect 367274 387922 367342 387978
rect 367398 387922 367494 387978
rect 366874 370350 367494 387922
rect 371648 382350 371968 382384
rect 371648 382294 371718 382350
rect 371774 382294 371842 382350
rect 371898 382294 371968 382350
rect 371648 382226 371968 382294
rect 371648 382170 371718 382226
rect 371774 382170 371842 382226
rect 371898 382170 371968 382226
rect 371648 382102 371968 382170
rect 371648 382046 371718 382102
rect 371774 382046 371842 382102
rect 371898 382046 371968 382102
rect 371648 381978 371968 382046
rect 371648 381922 371718 381978
rect 371774 381922 371842 381978
rect 371898 381922 371968 381978
rect 371648 381888 371968 381922
rect 381154 382350 381774 399922
rect 381154 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 381774 382350
rect 381154 382226 381774 382294
rect 381154 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 381774 382226
rect 381154 382102 381774 382170
rect 381154 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 381774 382102
rect 381154 381978 381774 382046
rect 381154 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 381774 381978
rect 366874 370294 366970 370350
rect 367026 370294 367094 370350
rect 367150 370294 367218 370350
rect 367274 370294 367342 370350
rect 367398 370294 367494 370350
rect 366874 370226 367494 370294
rect 366874 370170 366970 370226
rect 367026 370170 367094 370226
rect 367150 370170 367218 370226
rect 367274 370170 367342 370226
rect 367398 370170 367494 370226
rect 366874 370102 367494 370170
rect 366874 370046 366970 370102
rect 367026 370046 367094 370102
rect 367150 370046 367218 370102
rect 367274 370046 367342 370102
rect 367398 370046 367494 370102
rect 366874 369978 367494 370046
rect 366874 369922 366970 369978
rect 367026 369922 367094 369978
rect 367150 369922 367218 369978
rect 367274 369922 367342 369978
rect 367398 369922 367494 369978
rect 366874 352350 367494 369922
rect 371648 364350 371968 364384
rect 371648 364294 371718 364350
rect 371774 364294 371842 364350
rect 371898 364294 371968 364350
rect 371648 364226 371968 364294
rect 371648 364170 371718 364226
rect 371774 364170 371842 364226
rect 371898 364170 371968 364226
rect 371648 364102 371968 364170
rect 371648 364046 371718 364102
rect 371774 364046 371842 364102
rect 371898 364046 371968 364102
rect 371648 363978 371968 364046
rect 371648 363922 371718 363978
rect 371774 363922 371842 363978
rect 371898 363922 371968 363978
rect 371648 363888 371968 363922
rect 381154 364350 381774 381922
rect 381154 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 381774 364350
rect 381154 364226 381774 364294
rect 381154 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 381774 364226
rect 381154 364102 381774 364170
rect 381154 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 381774 364102
rect 381154 363978 381774 364046
rect 381154 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 381774 363978
rect 366874 352294 366970 352350
rect 367026 352294 367094 352350
rect 367150 352294 367218 352350
rect 367274 352294 367342 352350
rect 367398 352294 367494 352350
rect 366874 352226 367494 352294
rect 366874 352170 366970 352226
rect 367026 352170 367094 352226
rect 367150 352170 367218 352226
rect 367274 352170 367342 352226
rect 367398 352170 367494 352226
rect 366874 352102 367494 352170
rect 366874 352046 366970 352102
rect 367026 352046 367094 352102
rect 367150 352046 367218 352102
rect 367274 352046 367342 352102
rect 367398 352046 367494 352102
rect 366874 351978 367494 352046
rect 366874 351922 366970 351978
rect 367026 351922 367094 351978
rect 367150 351922 367218 351978
rect 367274 351922 367342 351978
rect 367398 351922 367494 351978
rect 366874 334350 367494 351922
rect 371648 346350 371968 346384
rect 371648 346294 371718 346350
rect 371774 346294 371842 346350
rect 371898 346294 371968 346350
rect 371648 346226 371968 346294
rect 371648 346170 371718 346226
rect 371774 346170 371842 346226
rect 371898 346170 371968 346226
rect 371648 346102 371968 346170
rect 371648 346046 371718 346102
rect 371774 346046 371842 346102
rect 371898 346046 371968 346102
rect 371648 345978 371968 346046
rect 371648 345922 371718 345978
rect 371774 345922 371842 345978
rect 371898 345922 371968 345978
rect 371648 345888 371968 345922
rect 381154 346350 381774 363922
rect 381154 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 381774 346350
rect 381154 346226 381774 346294
rect 381154 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 381774 346226
rect 381154 346102 381774 346170
rect 381154 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 381774 346102
rect 381154 345978 381774 346046
rect 381154 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 381774 345978
rect 366874 334294 366970 334350
rect 367026 334294 367094 334350
rect 367150 334294 367218 334350
rect 367274 334294 367342 334350
rect 367398 334294 367494 334350
rect 366874 334226 367494 334294
rect 366874 334170 366970 334226
rect 367026 334170 367094 334226
rect 367150 334170 367218 334226
rect 367274 334170 367342 334226
rect 367398 334170 367494 334226
rect 366874 334102 367494 334170
rect 366874 334046 366970 334102
rect 367026 334046 367094 334102
rect 367150 334046 367218 334102
rect 367274 334046 367342 334102
rect 367398 334046 367494 334102
rect 366874 333978 367494 334046
rect 366874 333922 366970 333978
rect 367026 333922 367094 333978
rect 367150 333922 367218 333978
rect 367274 333922 367342 333978
rect 367398 333922 367494 333978
rect 366874 316350 367494 333922
rect 371648 328350 371968 328384
rect 371648 328294 371718 328350
rect 371774 328294 371842 328350
rect 371898 328294 371968 328350
rect 371648 328226 371968 328294
rect 371648 328170 371718 328226
rect 371774 328170 371842 328226
rect 371898 328170 371968 328226
rect 371648 328102 371968 328170
rect 371648 328046 371718 328102
rect 371774 328046 371842 328102
rect 371898 328046 371968 328102
rect 371648 327978 371968 328046
rect 371648 327922 371718 327978
rect 371774 327922 371842 327978
rect 371898 327922 371968 327978
rect 371648 327888 371968 327922
rect 381154 328350 381774 345922
rect 381154 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 381774 328350
rect 381154 328226 381774 328294
rect 381154 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 381774 328226
rect 381154 328102 381774 328170
rect 381154 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 381774 328102
rect 381154 327978 381774 328046
rect 381154 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 381774 327978
rect 366874 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 367494 316350
rect 366874 316226 367494 316294
rect 366874 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 367494 316226
rect 366874 316102 367494 316170
rect 366874 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 367494 316102
rect 366874 315978 367494 316046
rect 366874 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 367494 315978
rect 366874 298350 367494 315922
rect 371648 310350 371968 310384
rect 371648 310294 371718 310350
rect 371774 310294 371842 310350
rect 371898 310294 371968 310350
rect 371648 310226 371968 310294
rect 371648 310170 371718 310226
rect 371774 310170 371842 310226
rect 371898 310170 371968 310226
rect 371648 310102 371968 310170
rect 371648 310046 371718 310102
rect 371774 310046 371842 310102
rect 371898 310046 371968 310102
rect 371648 309978 371968 310046
rect 371648 309922 371718 309978
rect 371774 309922 371842 309978
rect 371898 309922 371968 309978
rect 371648 309888 371968 309922
rect 381154 310350 381774 327922
rect 381154 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 381774 310350
rect 381154 310226 381774 310294
rect 381154 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 381774 310226
rect 381154 310102 381774 310170
rect 381154 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 381774 310102
rect 381154 309978 381774 310046
rect 381154 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 381774 309978
rect 366874 298294 366970 298350
rect 367026 298294 367094 298350
rect 367150 298294 367218 298350
rect 367274 298294 367342 298350
rect 367398 298294 367494 298350
rect 366874 298226 367494 298294
rect 366874 298170 366970 298226
rect 367026 298170 367094 298226
rect 367150 298170 367218 298226
rect 367274 298170 367342 298226
rect 367398 298170 367494 298226
rect 366874 298102 367494 298170
rect 366874 298046 366970 298102
rect 367026 298046 367094 298102
rect 367150 298046 367218 298102
rect 367274 298046 367342 298102
rect 367398 298046 367494 298102
rect 366874 297978 367494 298046
rect 366874 297922 366970 297978
rect 367026 297922 367094 297978
rect 367150 297922 367218 297978
rect 367274 297922 367342 297978
rect 367398 297922 367494 297978
rect 366874 280350 367494 297922
rect 371648 292350 371968 292384
rect 371648 292294 371718 292350
rect 371774 292294 371842 292350
rect 371898 292294 371968 292350
rect 371648 292226 371968 292294
rect 371648 292170 371718 292226
rect 371774 292170 371842 292226
rect 371898 292170 371968 292226
rect 371648 292102 371968 292170
rect 371648 292046 371718 292102
rect 371774 292046 371842 292102
rect 371898 292046 371968 292102
rect 371648 291978 371968 292046
rect 371648 291922 371718 291978
rect 371774 291922 371842 291978
rect 371898 291922 371968 291978
rect 371648 291888 371968 291922
rect 381154 292350 381774 309922
rect 381154 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 381774 292350
rect 381154 292226 381774 292294
rect 381154 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 381774 292226
rect 381154 292102 381774 292170
rect 381154 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 381774 292102
rect 381154 291978 381774 292046
rect 381154 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 381774 291978
rect 366874 280294 366970 280350
rect 367026 280294 367094 280350
rect 367150 280294 367218 280350
rect 367274 280294 367342 280350
rect 367398 280294 367494 280350
rect 366874 280226 367494 280294
rect 366874 280170 366970 280226
rect 367026 280170 367094 280226
rect 367150 280170 367218 280226
rect 367274 280170 367342 280226
rect 367398 280170 367494 280226
rect 366874 280102 367494 280170
rect 366874 280046 366970 280102
rect 367026 280046 367094 280102
rect 367150 280046 367218 280102
rect 367274 280046 367342 280102
rect 367398 280046 367494 280102
rect 366874 279978 367494 280046
rect 366874 279922 366970 279978
rect 367026 279922 367094 279978
rect 367150 279922 367218 279978
rect 367274 279922 367342 279978
rect 367398 279922 367494 279978
rect 366874 262350 367494 279922
rect 371648 274350 371968 274384
rect 371648 274294 371718 274350
rect 371774 274294 371842 274350
rect 371898 274294 371968 274350
rect 371648 274226 371968 274294
rect 371648 274170 371718 274226
rect 371774 274170 371842 274226
rect 371898 274170 371968 274226
rect 371648 274102 371968 274170
rect 371648 274046 371718 274102
rect 371774 274046 371842 274102
rect 371898 274046 371968 274102
rect 371648 273978 371968 274046
rect 371648 273922 371718 273978
rect 371774 273922 371842 273978
rect 371898 273922 371968 273978
rect 371648 273888 371968 273922
rect 381154 274350 381774 291922
rect 381154 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 381774 274350
rect 381154 274226 381774 274294
rect 381154 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 381774 274226
rect 381154 274102 381774 274170
rect 381154 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 381774 274102
rect 381154 273978 381774 274046
rect 381154 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 381774 273978
rect 366874 262294 366970 262350
rect 367026 262294 367094 262350
rect 367150 262294 367218 262350
rect 367274 262294 367342 262350
rect 367398 262294 367494 262350
rect 366874 262226 367494 262294
rect 366874 262170 366970 262226
rect 367026 262170 367094 262226
rect 367150 262170 367218 262226
rect 367274 262170 367342 262226
rect 367398 262170 367494 262226
rect 366874 262102 367494 262170
rect 366874 262046 366970 262102
rect 367026 262046 367094 262102
rect 367150 262046 367218 262102
rect 367274 262046 367342 262102
rect 367398 262046 367494 262102
rect 366874 261978 367494 262046
rect 366874 261922 366970 261978
rect 367026 261922 367094 261978
rect 367150 261922 367218 261978
rect 367274 261922 367342 261978
rect 367398 261922 367494 261978
rect 366874 244350 367494 261922
rect 371648 256350 371968 256384
rect 371648 256294 371718 256350
rect 371774 256294 371842 256350
rect 371898 256294 371968 256350
rect 371648 256226 371968 256294
rect 371648 256170 371718 256226
rect 371774 256170 371842 256226
rect 371898 256170 371968 256226
rect 371648 256102 371968 256170
rect 371648 256046 371718 256102
rect 371774 256046 371842 256102
rect 371898 256046 371968 256102
rect 371648 255978 371968 256046
rect 371648 255922 371718 255978
rect 371774 255922 371842 255978
rect 371898 255922 371968 255978
rect 371648 255888 371968 255922
rect 381154 256350 381774 273922
rect 381154 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 381774 256350
rect 381154 256226 381774 256294
rect 381154 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 381774 256226
rect 381154 256102 381774 256170
rect 381154 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 381774 256102
rect 381154 255978 381774 256046
rect 381154 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 381774 255978
rect 366874 244294 366970 244350
rect 367026 244294 367094 244350
rect 367150 244294 367218 244350
rect 367274 244294 367342 244350
rect 367398 244294 367494 244350
rect 366874 244226 367494 244294
rect 366874 244170 366970 244226
rect 367026 244170 367094 244226
rect 367150 244170 367218 244226
rect 367274 244170 367342 244226
rect 367398 244170 367494 244226
rect 366874 244102 367494 244170
rect 366874 244046 366970 244102
rect 367026 244046 367094 244102
rect 367150 244046 367218 244102
rect 367274 244046 367342 244102
rect 367398 244046 367494 244102
rect 366874 243978 367494 244046
rect 366874 243922 366970 243978
rect 367026 243922 367094 243978
rect 367150 243922 367218 243978
rect 367274 243922 367342 243978
rect 367398 243922 367494 243978
rect 366874 226350 367494 243922
rect 371648 238350 371968 238384
rect 371648 238294 371718 238350
rect 371774 238294 371842 238350
rect 371898 238294 371968 238350
rect 371648 238226 371968 238294
rect 371648 238170 371718 238226
rect 371774 238170 371842 238226
rect 371898 238170 371968 238226
rect 371648 238102 371968 238170
rect 371648 238046 371718 238102
rect 371774 238046 371842 238102
rect 371898 238046 371968 238102
rect 371648 237978 371968 238046
rect 371648 237922 371718 237978
rect 371774 237922 371842 237978
rect 371898 237922 371968 237978
rect 371648 237888 371968 237922
rect 381154 238350 381774 255922
rect 381154 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 381774 238350
rect 381154 238226 381774 238294
rect 381154 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 381774 238226
rect 381154 238102 381774 238170
rect 381154 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 381774 238102
rect 381154 237978 381774 238046
rect 381154 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 381774 237978
rect 366874 226294 366970 226350
rect 367026 226294 367094 226350
rect 367150 226294 367218 226350
rect 367274 226294 367342 226350
rect 367398 226294 367494 226350
rect 366874 226226 367494 226294
rect 366874 226170 366970 226226
rect 367026 226170 367094 226226
rect 367150 226170 367218 226226
rect 367274 226170 367342 226226
rect 367398 226170 367494 226226
rect 366874 226102 367494 226170
rect 366874 226046 366970 226102
rect 367026 226046 367094 226102
rect 367150 226046 367218 226102
rect 367274 226046 367342 226102
rect 367398 226046 367494 226102
rect 366874 225978 367494 226046
rect 366874 225922 366970 225978
rect 367026 225922 367094 225978
rect 367150 225922 367218 225978
rect 367274 225922 367342 225978
rect 367398 225922 367494 225978
rect 366874 208350 367494 225922
rect 371648 220350 371968 220384
rect 371648 220294 371718 220350
rect 371774 220294 371842 220350
rect 371898 220294 371968 220350
rect 371648 220226 371968 220294
rect 371648 220170 371718 220226
rect 371774 220170 371842 220226
rect 371898 220170 371968 220226
rect 371648 220102 371968 220170
rect 371648 220046 371718 220102
rect 371774 220046 371842 220102
rect 371898 220046 371968 220102
rect 371648 219978 371968 220046
rect 371648 219922 371718 219978
rect 371774 219922 371842 219978
rect 371898 219922 371968 219978
rect 371648 219888 371968 219922
rect 381154 220350 381774 237922
rect 381154 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 381774 220350
rect 381154 220226 381774 220294
rect 381154 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 381774 220226
rect 381154 220102 381774 220170
rect 381154 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 381774 220102
rect 381154 219978 381774 220046
rect 381154 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 381774 219978
rect 366874 208294 366970 208350
rect 367026 208294 367094 208350
rect 367150 208294 367218 208350
rect 367274 208294 367342 208350
rect 367398 208294 367494 208350
rect 366874 208226 367494 208294
rect 366874 208170 366970 208226
rect 367026 208170 367094 208226
rect 367150 208170 367218 208226
rect 367274 208170 367342 208226
rect 367398 208170 367494 208226
rect 366874 208102 367494 208170
rect 366874 208046 366970 208102
rect 367026 208046 367094 208102
rect 367150 208046 367218 208102
rect 367274 208046 367342 208102
rect 367398 208046 367494 208102
rect 366874 207978 367494 208046
rect 366874 207922 366970 207978
rect 367026 207922 367094 207978
rect 367150 207922 367218 207978
rect 367274 207922 367342 207978
rect 367398 207922 367494 207978
rect 366874 190350 367494 207922
rect 371648 202350 371968 202384
rect 371648 202294 371718 202350
rect 371774 202294 371842 202350
rect 371898 202294 371968 202350
rect 371648 202226 371968 202294
rect 371648 202170 371718 202226
rect 371774 202170 371842 202226
rect 371898 202170 371968 202226
rect 371648 202102 371968 202170
rect 371648 202046 371718 202102
rect 371774 202046 371842 202102
rect 371898 202046 371968 202102
rect 371648 201978 371968 202046
rect 371648 201922 371718 201978
rect 371774 201922 371842 201978
rect 371898 201922 371968 201978
rect 371648 201888 371968 201922
rect 381154 202350 381774 219922
rect 381154 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 381774 202350
rect 381154 202226 381774 202294
rect 381154 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 381774 202226
rect 381154 202102 381774 202170
rect 381154 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 381774 202102
rect 381154 201978 381774 202046
rect 381154 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 381774 201978
rect 366874 190294 366970 190350
rect 367026 190294 367094 190350
rect 367150 190294 367218 190350
rect 367274 190294 367342 190350
rect 367398 190294 367494 190350
rect 366874 190226 367494 190294
rect 366874 190170 366970 190226
rect 367026 190170 367094 190226
rect 367150 190170 367218 190226
rect 367274 190170 367342 190226
rect 367398 190170 367494 190226
rect 366874 190102 367494 190170
rect 366874 190046 366970 190102
rect 367026 190046 367094 190102
rect 367150 190046 367218 190102
rect 367274 190046 367342 190102
rect 367398 190046 367494 190102
rect 366874 189978 367494 190046
rect 366874 189922 366970 189978
rect 367026 189922 367094 189978
rect 367150 189922 367218 189978
rect 367274 189922 367342 189978
rect 367398 189922 367494 189978
rect 366874 172350 367494 189922
rect 371648 184350 371968 184384
rect 371648 184294 371718 184350
rect 371774 184294 371842 184350
rect 371898 184294 371968 184350
rect 371648 184226 371968 184294
rect 371648 184170 371718 184226
rect 371774 184170 371842 184226
rect 371898 184170 371968 184226
rect 371648 184102 371968 184170
rect 371648 184046 371718 184102
rect 371774 184046 371842 184102
rect 371898 184046 371968 184102
rect 371648 183978 371968 184046
rect 371648 183922 371718 183978
rect 371774 183922 371842 183978
rect 371898 183922 371968 183978
rect 371648 183888 371968 183922
rect 381154 184350 381774 201922
rect 381154 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 381774 184350
rect 381154 184226 381774 184294
rect 381154 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 381774 184226
rect 381154 184102 381774 184170
rect 381154 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 381774 184102
rect 381154 183978 381774 184046
rect 381154 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 381774 183978
rect 366874 172294 366970 172350
rect 367026 172294 367094 172350
rect 367150 172294 367218 172350
rect 367274 172294 367342 172350
rect 367398 172294 367494 172350
rect 366874 172226 367494 172294
rect 366874 172170 366970 172226
rect 367026 172170 367094 172226
rect 367150 172170 367218 172226
rect 367274 172170 367342 172226
rect 367398 172170 367494 172226
rect 366874 172102 367494 172170
rect 366874 172046 366970 172102
rect 367026 172046 367094 172102
rect 367150 172046 367218 172102
rect 367274 172046 367342 172102
rect 367398 172046 367494 172102
rect 366874 171978 367494 172046
rect 366874 171922 366970 171978
rect 367026 171922 367094 171978
rect 367150 171922 367218 171978
rect 367274 171922 367342 171978
rect 367398 171922 367494 171978
rect 366874 154350 367494 171922
rect 371648 166350 371968 166384
rect 371648 166294 371718 166350
rect 371774 166294 371842 166350
rect 371898 166294 371968 166350
rect 371648 166226 371968 166294
rect 371648 166170 371718 166226
rect 371774 166170 371842 166226
rect 371898 166170 371968 166226
rect 371648 166102 371968 166170
rect 371648 166046 371718 166102
rect 371774 166046 371842 166102
rect 371898 166046 371968 166102
rect 371648 165978 371968 166046
rect 371648 165922 371718 165978
rect 371774 165922 371842 165978
rect 371898 165922 371968 165978
rect 371648 165888 371968 165922
rect 381154 166350 381774 183922
rect 381154 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 381774 166350
rect 381154 166226 381774 166294
rect 381154 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 381774 166226
rect 381154 166102 381774 166170
rect 381154 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 381774 166102
rect 381154 165978 381774 166046
rect 381154 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 381774 165978
rect 366874 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 367494 154350
rect 366874 154226 367494 154294
rect 366874 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 367494 154226
rect 366874 154102 367494 154170
rect 366874 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 367494 154102
rect 366874 153978 367494 154046
rect 366874 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 367494 153978
rect 366874 136350 367494 153922
rect 371648 148350 371968 148384
rect 371648 148294 371718 148350
rect 371774 148294 371842 148350
rect 371898 148294 371968 148350
rect 371648 148226 371968 148294
rect 371648 148170 371718 148226
rect 371774 148170 371842 148226
rect 371898 148170 371968 148226
rect 371648 148102 371968 148170
rect 371648 148046 371718 148102
rect 371774 148046 371842 148102
rect 371898 148046 371968 148102
rect 371648 147978 371968 148046
rect 371648 147922 371718 147978
rect 371774 147922 371842 147978
rect 371898 147922 371968 147978
rect 371648 147888 371968 147922
rect 381154 148350 381774 165922
rect 381154 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 381774 148350
rect 381154 148226 381774 148294
rect 381154 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 381774 148226
rect 381154 148102 381774 148170
rect 381154 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 381774 148102
rect 381154 147978 381774 148046
rect 381154 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 381774 147978
rect 366874 136294 366970 136350
rect 367026 136294 367094 136350
rect 367150 136294 367218 136350
rect 367274 136294 367342 136350
rect 367398 136294 367494 136350
rect 366874 136226 367494 136294
rect 366874 136170 366970 136226
rect 367026 136170 367094 136226
rect 367150 136170 367218 136226
rect 367274 136170 367342 136226
rect 367398 136170 367494 136226
rect 366874 136102 367494 136170
rect 366874 136046 366970 136102
rect 367026 136046 367094 136102
rect 367150 136046 367218 136102
rect 367274 136046 367342 136102
rect 367398 136046 367494 136102
rect 366874 135978 367494 136046
rect 366874 135922 366970 135978
rect 367026 135922 367094 135978
rect 367150 135922 367218 135978
rect 367274 135922 367342 135978
rect 367398 135922 367494 135978
rect 366874 118350 367494 135922
rect 371648 130350 371968 130384
rect 371648 130294 371718 130350
rect 371774 130294 371842 130350
rect 371898 130294 371968 130350
rect 371648 130226 371968 130294
rect 371648 130170 371718 130226
rect 371774 130170 371842 130226
rect 371898 130170 371968 130226
rect 371648 130102 371968 130170
rect 371648 130046 371718 130102
rect 371774 130046 371842 130102
rect 371898 130046 371968 130102
rect 371648 129978 371968 130046
rect 371648 129922 371718 129978
rect 371774 129922 371842 129978
rect 371898 129922 371968 129978
rect 371648 129888 371968 129922
rect 381154 130350 381774 147922
rect 381154 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 381774 130350
rect 381154 130226 381774 130294
rect 381154 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 381774 130226
rect 381154 130102 381774 130170
rect 381154 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 381774 130102
rect 381154 129978 381774 130046
rect 381154 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 381774 129978
rect 366874 118294 366970 118350
rect 367026 118294 367094 118350
rect 367150 118294 367218 118350
rect 367274 118294 367342 118350
rect 367398 118294 367494 118350
rect 366874 118226 367494 118294
rect 366874 118170 366970 118226
rect 367026 118170 367094 118226
rect 367150 118170 367218 118226
rect 367274 118170 367342 118226
rect 367398 118170 367494 118226
rect 366874 118102 367494 118170
rect 366874 118046 366970 118102
rect 367026 118046 367094 118102
rect 367150 118046 367218 118102
rect 367274 118046 367342 118102
rect 367398 118046 367494 118102
rect 366874 117978 367494 118046
rect 366874 117922 366970 117978
rect 367026 117922 367094 117978
rect 367150 117922 367218 117978
rect 367274 117922 367342 117978
rect 367398 117922 367494 117978
rect 366874 100350 367494 117922
rect 371648 112350 371968 112384
rect 371648 112294 371718 112350
rect 371774 112294 371842 112350
rect 371898 112294 371968 112350
rect 371648 112226 371968 112294
rect 371648 112170 371718 112226
rect 371774 112170 371842 112226
rect 371898 112170 371968 112226
rect 371648 112102 371968 112170
rect 371648 112046 371718 112102
rect 371774 112046 371842 112102
rect 371898 112046 371968 112102
rect 371648 111978 371968 112046
rect 371648 111922 371718 111978
rect 371774 111922 371842 111978
rect 371898 111922 371968 111978
rect 371648 111888 371968 111922
rect 381154 112350 381774 129922
rect 381154 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 381774 112350
rect 381154 112226 381774 112294
rect 381154 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 381774 112226
rect 381154 112102 381774 112170
rect 381154 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 381774 112102
rect 381154 111978 381774 112046
rect 381154 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 381774 111978
rect 366874 100294 366970 100350
rect 367026 100294 367094 100350
rect 367150 100294 367218 100350
rect 367274 100294 367342 100350
rect 367398 100294 367494 100350
rect 366874 100226 367494 100294
rect 366874 100170 366970 100226
rect 367026 100170 367094 100226
rect 367150 100170 367218 100226
rect 367274 100170 367342 100226
rect 367398 100170 367494 100226
rect 366874 100102 367494 100170
rect 366874 100046 366970 100102
rect 367026 100046 367094 100102
rect 367150 100046 367218 100102
rect 367274 100046 367342 100102
rect 367398 100046 367494 100102
rect 366874 99978 367494 100046
rect 366874 99922 366970 99978
rect 367026 99922 367094 99978
rect 367150 99922 367218 99978
rect 367274 99922 367342 99978
rect 367398 99922 367494 99978
rect 366874 82350 367494 99922
rect 371648 94350 371968 94384
rect 371648 94294 371718 94350
rect 371774 94294 371842 94350
rect 371898 94294 371968 94350
rect 371648 94226 371968 94294
rect 371648 94170 371718 94226
rect 371774 94170 371842 94226
rect 371898 94170 371968 94226
rect 371648 94102 371968 94170
rect 371648 94046 371718 94102
rect 371774 94046 371842 94102
rect 371898 94046 371968 94102
rect 371648 93978 371968 94046
rect 371648 93922 371718 93978
rect 371774 93922 371842 93978
rect 371898 93922 371968 93978
rect 371648 93888 371968 93922
rect 381154 94350 381774 111922
rect 381154 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 381774 94350
rect 381154 94226 381774 94294
rect 381154 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 381774 94226
rect 381154 94102 381774 94170
rect 381154 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 381774 94102
rect 381154 93978 381774 94046
rect 381154 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 381774 93978
rect 366874 82294 366970 82350
rect 367026 82294 367094 82350
rect 367150 82294 367218 82350
rect 367274 82294 367342 82350
rect 367398 82294 367494 82350
rect 366874 82226 367494 82294
rect 366874 82170 366970 82226
rect 367026 82170 367094 82226
rect 367150 82170 367218 82226
rect 367274 82170 367342 82226
rect 367398 82170 367494 82226
rect 366874 82102 367494 82170
rect 366874 82046 366970 82102
rect 367026 82046 367094 82102
rect 367150 82046 367218 82102
rect 367274 82046 367342 82102
rect 367398 82046 367494 82102
rect 366874 81978 367494 82046
rect 366874 81922 366970 81978
rect 367026 81922 367094 81978
rect 367150 81922 367218 81978
rect 367274 81922 367342 81978
rect 367398 81922 367494 81978
rect 366874 64350 367494 81922
rect 371648 76350 371968 76384
rect 371648 76294 371718 76350
rect 371774 76294 371842 76350
rect 371898 76294 371968 76350
rect 371648 76226 371968 76294
rect 371648 76170 371718 76226
rect 371774 76170 371842 76226
rect 371898 76170 371968 76226
rect 371648 76102 371968 76170
rect 371648 76046 371718 76102
rect 371774 76046 371842 76102
rect 371898 76046 371968 76102
rect 371648 75978 371968 76046
rect 371648 75922 371718 75978
rect 371774 75922 371842 75978
rect 371898 75922 371968 75978
rect 371648 75888 371968 75922
rect 381154 76350 381774 93922
rect 381154 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 381774 76350
rect 381154 76226 381774 76294
rect 381154 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 381774 76226
rect 381154 76102 381774 76170
rect 381154 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 381774 76102
rect 381154 75978 381774 76046
rect 381154 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 381774 75978
rect 366874 64294 366970 64350
rect 367026 64294 367094 64350
rect 367150 64294 367218 64350
rect 367274 64294 367342 64350
rect 367398 64294 367494 64350
rect 366874 64226 367494 64294
rect 366874 64170 366970 64226
rect 367026 64170 367094 64226
rect 367150 64170 367218 64226
rect 367274 64170 367342 64226
rect 367398 64170 367494 64226
rect 366874 64102 367494 64170
rect 366874 64046 366970 64102
rect 367026 64046 367094 64102
rect 367150 64046 367218 64102
rect 367274 64046 367342 64102
rect 367398 64046 367494 64102
rect 366874 63978 367494 64046
rect 366874 63922 366970 63978
rect 367026 63922 367094 63978
rect 367150 63922 367218 63978
rect 367274 63922 367342 63978
rect 367398 63922 367494 63978
rect 366874 46350 367494 63922
rect 366874 46294 366970 46350
rect 367026 46294 367094 46350
rect 367150 46294 367218 46350
rect 367274 46294 367342 46350
rect 367398 46294 367494 46350
rect 366874 46226 367494 46294
rect 366874 46170 366970 46226
rect 367026 46170 367094 46226
rect 367150 46170 367218 46226
rect 367274 46170 367342 46226
rect 367398 46170 367494 46226
rect 366874 46102 367494 46170
rect 366874 46046 366970 46102
rect 367026 46046 367094 46102
rect 367150 46046 367218 46102
rect 367274 46046 367342 46102
rect 367398 46046 367494 46102
rect 366874 45978 367494 46046
rect 366874 45922 366970 45978
rect 367026 45922 367094 45978
rect 367150 45922 367218 45978
rect 367274 45922 367342 45978
rect 367398 45922 367494 45978
rect 366874 28350 367494 45922
rect 366874 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 367494 28350
rect 366874 28226 367494 28294
rect 366874 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 367494 28226
rect 366874 28102 367494 28170
rect 366874 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 367494 28102
rect 366874 27978 367494 28046
rect 366874 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 367494 27978
rect 366874 10350 367494 27922
rect 366874 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 367494 10350
rect 366874 10226 367494 10294
rect 366874 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 367494 10226
rect 366874 10102 367494 10170
rect 366874 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 367494 10102
rect 366874 9978 367494 10046
rect 366874 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 367494 9978
rect 366874 -1120 367494 9922
rect 366874 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 367494 -1120
rect 366874 -1244 367494 -1176
rect 366874 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 367494 -1244
rect 366874 -1368 367494 -1300
rect 366874 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 367494 -1368
rect 366874 -1492 367494 -1424
rect 366874 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 367494 -1492
rect 366874 -1644 367494 -1548
rect 381154 58350 381774 75922
rect 381154 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 381774 58350
rect 381154 58226 381774 58294
rect 381154 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 381774 58226
rect 381154 58102 381774 58170
rect 381154 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 381774 58102
rect 381154 57978 381774 58046
rect 381154 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 381774 57978
rect 381154 40350 381774 57922
rect 381154 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 381774 40350
rect 381154 40226 381774 40294
rect 381154 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 381774 40226
rect 381154 40102 381774 40170
rect 381154 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 381774 40102
rect 381154 39978 381774 40046
rect 381154 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 381774 39978
rect 381154 22350 381774 39922
rect 381154 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 381774 22350
rect 381154 22226 381774 22294
rect 381154 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 381774 22226
rect 381154 22102 381774 22170
rect 381154 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 381774 22102
rect 381154 21978 381774 22046
rect 381154 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 381774 21978
rect 381154 4350 381774 21922
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 598172 385494 598268
rect 384874 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 385494 598172
rect 384874 598048 385494 598116
rect 384874 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 385494 598048
rect 384874 597924 385494 597992
rect 384874 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 385494 597924
rect 384874 597800 385494 597868
rect 384874 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 385494 597800
rect 384874 586350 385494 597744
rect 384874 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 385494 586350
rect 384874 586226 385494 586294
rect 384874 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 385494 586226
rect 384874 586102 385494 586170
rect 384874 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 385494 586102
rect 384874 585978 385494 586046
rect 384874 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 385494 585978
rect 384874 568350 385494 585922
rect 384874 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 385494 568350
rect 384874 568226 385494 568294
rect 384874 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 385494 568226
rect 384874 568102 385494 568170
rect 384874 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 385494 568102
rect 384874 567978 385494 568046
rect 384874 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 385494 567978
rect 384874 550350 385494 567922
rect 384874 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 385494 550350
rect 384874 550226 385494 550294
rect 384874 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 385494 550226
rect 384874 550102 385494 550170
rect 384874 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 385494 550102
rect 384874 549978 385494 550046
rect 384874 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 385494 549978
rect 384874 532350 385494 549922
rect 384874 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 385494 532350
rect 384874 532226 385494 532294
rect 384874 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 385494 532226
rect 384874 532102 385494 532170
rect 384874 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 385494 532102
rect 384874 531978 385494 532046
rect 384874 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 385494 531978
rect 384874 514350 385494 531922
rect 384874 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 385494 514350
rect 384874 514226 385494 514294
rect 384874 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 385494 514226
rect 384874 514102 385494 514170
rect 384874 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 385494 514102
rect 384874 513978 385494 514046
rect 384874 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 385494 513978
rect 384874 496350 385494 513922
rect 384874 496294 384970 496350
rect 385026 496294 385094 496350
rect 385150 496294 385218 496350
rect 385274 496294 385342 496350
rect 385398 496294 385494 496350
rect 384874 496226 385494 496294
rect 384874 496170 384970 496226
rect 385026 496170 385094 496226
rect 385150 496170 385218 496226
rect 385274 496170 385342 496226
rect 385398 496170 385494 496226
rect 384874 496102 385494 496170
rect 384874 496046 384970 496102
rect 385026 496046 385094 496102
rect 385150 496046 385218 496102
rect 385274 496046 385342 496102
rect 385398 496046 385494 496102
rect 384874 495978 385494 496046
rect 384874 495922 384970 495978
rect 385026 495922 385094 495978
rect 385150 495922 385218 495978
rect 385274 495922 385342 495978
rect 385398 495922 385494 495978
rect 384874 478350 385494 495922
rect 384874 478294 384970 478350
rect 385026 478294 385094 478350
rect 385150 478294 385218 478350
rect 385274 478294 385342 478350
rect 385398 478294 385494 478350
rect 384874 478226 385494 478294
rect 384874 478170 384970 478226
rect 385026 478170 385094 478226
rect 385150 478170 385218 478226
rect 385274 478170 385342 478226
rect 385398 478170 385494 478226
rect 384874 478102 385494 478170
rect 384874 478046 384970 478102
rect 385026 478046 385094 478102
rect 385150 478046 385218 478102
rect 385274 478046 385342 478102
rect 385398 478046 385494 478102
rect 384874 477978 385494 478046
rect 384874 477922 384970 477978
rect 385026 477922 385094 477978
rect 385150 477922 385218 477978
rect 385274 477922 385342 477978
rect 385398 477922 385494 477978
rect 384874 460350 385494 477922
rect 384874 460294 384970 460350
rect 385026 460294 385094 460350
rect 385150 460294 385218 460350
rect 385274 460294 385342 460350
rect 385398 460294 385494 460350
rect 384874 460226 385494 460294
rect 384874 460170 384970 460226
rect 385026 460170 385094 460226
rect 385150 460170 385218 460226
rect 385274 460170 385342 460226
rect 385398 460170 385494 460226
rect 384874 460102 385494 460170
rect 384874 460046 384970 460102
rect 385026 460046 385094 460102
rect 385150 460046 385218 460102
rect 385274 460046 385342 460102
rect 385398 460046 385494 460102
rect 384874 459978 385494 460046
rect 384874 459922 384970 459978
rect 385026 459922 385094 459978
rect 385150 459922 385218 459978
rect 385274 459922 385342 459978
rect 385398 459922 385494 459978
rect 384874 442350 385494 459922
rect 384874 442294 384970 442350
rect 385026 442294 385094 442350
rect 385150 442294 385218 442350
rect 385274 442294 385342 442350
rect 385398 442294 385494 442350
rect 384874 442226 385494 442294
rect 384874 442170 384970 442226
rect 385026 442170 385094 442226
rect 385150 442170 385218 442226
rect 385274 442170 385342 442226
rect 385398 442170 385494 442226
rect 384874 442102 385494 442170
rect 384874 442046 384970 442102
rect 385026 442046 385094 442102
rect 385150 442046 385218 442102
rect 385274 442046 385342 442102
rect 385398 442046 385494 442102
rect 384874 441978 385494 442046
rect 384874 441922 384970 441978
rect 385026 441922 385094 441978
rect 385150 441922 385218 441978
rect 385274 441922 385342 441978
rect 385398 441922 385494 441978
rect 384874 424350 385494 441922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 526350 399774 543922
rect 399154 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 399774 526350
rect 399154 526226 399774 526294
rect 399154 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 399774 526226
rect 399154 526102 399774 526170
rect 399154 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 399774 526102
rect 399154 525978 399774 526046
rect 399154 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 399774 525978
rect 399154 508350 399774 525922
rect 399154 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 399774 508350
rect 399154 508226 399774 508294
rect 399154 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 399774 508226
rect 399154 508102 399774 508170
rect 399154 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 399774 508102
rect 399154 507978 399774 508046
rect 399154 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 399774 507978
rect 399154 490350 399774 507922
rect 399154 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 399774 490350
rect 399154 490226 399774 490294
rect 399154 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 399774 490226
rect 399154 490102 399774 490170
rect 399154 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 399774 490102
rect 399154 489978 399774 490046
rect 399154 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 399774 489978
rect 399154 472350 399774 489922
rect 399154 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 399774 472350
rect 399154 472226 399774 472294
rect 399154 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 399774 472226
rect 399154 472102 399774 472170
rect 399154 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 399774 472102
rect 399154 471978 399774 472046
rect 399154 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 399774 471978
rect 399154 454350 399774 471922
rect 399154 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 399774 454350
rect 399154 454226 399774 454294
rect 399154 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 399774 454226
rect 399154 454102 399774 454170
rect 399154 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 399774 454102
rect 399154 453978 399774 454046
rect 399154 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 399774 453978
rect 399154 436350 399774 453922
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 514350 403494 531922
rect 402874 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 403494 514350
rect 402874 514226 403494 514294
rect 402874 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 403494 514226
rect 402874 514102 403494 514170
rect 402874 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 403494 514102
rect 402874 513978 403494 514046
rect 402874 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 403494 513978
rect 402874 496350 403494 513922
rect 402874 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 403494 496350
rect 402874 496226 403494 496294
rect 402874 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 403494 496226
rect 402874 496102 403494 496170
rect 402874 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 403494 496102
rect 402874 495978 403494 496046
rect 402874 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 403494 495978
rect 402874 478350 403494 495922
rect 402874 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 403494 478350
rect 402874 478226 403494 478294
rect 402874 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 403494 478226
rect 402874 478102 403494 478170
rect 402874 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 403494 478102
rect 402874 477978 403494 478046
rect 402874 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 403494 477978
rect 402874 460350 403494 477922
rect 402874 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 403494 460350
rect 402874 460226 403494 460294
rect 402874 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 403494 460226
rect 402874 460102 403494 460170
rect 402874 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 403494 460102
rect 402874 459978 403494 460046
rect 402874 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 403494 459978
rect 402874 442350 403494 459922
rect 402874 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 403494 442350
rect 402874 442226 403494 442294
rect 402874 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 403494 442226
rect 402874 442102 403494 442170
rect 402874 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 403494 442102
rect 402874 441978 403494 442046
rect 402874 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 403494 441978
rect 399154 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436294 399774 436350
rect 399154 436226 399774 436294
rect 399154 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436170 399774 436226
rect 399154 436102 399774 436170
rect 399154 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436046 399774 436102
rect 399154 435978 399774 436046
rect 399154 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435922 399774 435978
rect 384874 424294 384970 424350
rect 385026 424294 385094 424350
rect 385150 424294 385218 424350
rect 385274 424294 385342 424350
rect 385398 424294 385494 424350
rect 384874 424226 385494 424294
rect 384874 424170 384970 424226
rect 385026 424170 385094 424226
rect 385150 424170 385218 424226
rect 385274 424170 385342 424226
rect 385398 424170 385494 424226
rect 384874 424102 385494 424170
rect 384874 424046 384970 424102
rect 385026 424046 385094 424102
rect 385150 424046 385218 424102
rect 385274 424046 385342 424102
rect 385398 424046 385494 424102
rect 384874 423978 385494 424046
rect 384874 423922 384970 423978
rect 385026 423922 385094 423978
rect 385150 423922 385218 423978
rect 385274 423922 385342 423978
rect 385398 423922 385494 423978
rect 384874 406350 385494 423922
rect 387008 424350 387328 424384
rect 387008 424294 387078 424350
rect 387134 424294 387202 424350
rect 387258 424294 387328 424350
rect 387008 424226 387328 424294
rect 387008 424170 387078 424226
rect 387134 424170 387202 424226
rect 387258 424170 387328 424226
rect 387008 424102 387328 424170
rect 387008 424046 387078 424102
rect 387134 424046 387202 424102
rect 387258 424046 387328 424102
rect 387008 423978 387328 424046
rect 387008 423922 387078 423978
rect 387134 423922 387202 423978
rect 387258 423922 387328 423978
rect 387008 423888 387328 423922
rect 399154 418350 399774 435922
rect 402368 436317 402688 436380
rect 402368 436261 402438 436317
rect 402494 436261 402562 436317
rect 402618 436261 402688 436317
rect 402368 436193 402688 436261
rect 402368 436137 402438 436193
rect 402494 436137 402562 436193
rect 402618 436137 402688 436193
rect 402368 436069 402688 436137
rect 402368 436013 402438 436069
rect 402494 436013 402562 436069
rect 402618 436013 402688 436069
rect 402368 435945 402688 436013
rect 402368 435889 402438 435945
rect 402494 435889 402562 435945
rect 402618 435889 402688 435945
rect 402368 435826 402688 435889
rect 402874 424350 403494 441922
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 526350 417774 543922
rect 417154 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 417774 526350
rect 417154 526226 417774 526294
rect 417154 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 417774 526226
rect 417154 526102 417774 526170
rect 417154 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 417774 526102
rect 417154 525978 417774 526046
rect 417154 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 417774 525978
rect 417154 508350 417774 525922
rect 417154 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 417774 508350
rect 417154 508226 417774 508294
rect 417154 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 417774 508226
rect 417154 508102 417774 508170
rect 417154 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 417774 508102
rect 417154 507978 417774 508046
rect 417154 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 417774 507978
rect 417154 490350 417774 507922
rect 417154 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 417774 490350
rect 417154 490226 417774 490294
rect 417154 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 417774 490226
rect 417154 490102 417774 490170
rect 417154 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 417774 490102
rect 417154 489978 417774 490046
rect 417154 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 417774 489978
rect 417154 472350 417774 489922
rect 417154 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 417774 472350
rect 417154 472226 417774 472294
rect 417154 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 417774 472226
rect 417154 472102 417774 472170
rect 417154 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 417774 472102
rect 417154 471978 417774 472046
rect 417154 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 417774 471978
rect 417154 454350 417774 471922
rect 417154 454294 417250 454350
rect 417306 454294 417374 454350
rect 417430 454294 417498 454350
rect 417554 454294 417622 454350
rect 417678 454294 417774 454350
rect 417154 454226 417774 454294
rect 417154 454170 417250 454226
rect 417306 454170 417374 454226
rect 417430 454170 417498 454226
rect 417554 454170 417622 454226
rect 417678 454170 417774 454226
rect 417154 454102 417774 454170
rect 417154 454046 417250 454102
rect 417306 454046 417374 454102
rect 417430 454046 417498 454102
rect 417554 454046 417622 454102
rect 417678 454046 417774 454102
rect 417154 453978 417774 454046
rect 417154 453922 417250 453978
rect 417306 453922 417374 453978
rect 417430 453922 417498 453978
rect 417554 453922 417622 453978
rect 417678 453922 417774 453978
rect 417154 438436 417774 453922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 514350 421494 531922
rect 420874 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 421494 514350
rect 420874 514226 421494 514294
rect 420874 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 421494 514226
rect 420874 514102 421494 514170
rect 420874 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 421494 514102
rect 420874 513978 421494 514046
rect 420874 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 421494 513978
rect 420874 496350 421494 513922
rect 420874 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 421494 496350
rect 420874 496226 421494 496294
rect 420874 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 421494 496226
rect 420874 496102 421494 496170
rect 420874 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 421494 496102
rect 420874 495978 421494 496046
rect 420874 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 421494 495978
rect 420874 478350 421494 495922
rect 420874 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 421494 478350
rect 420874 478226 421494 478294
rect 420874 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 421494 478226
rect 420874 478102 421494 478170
rect 420874 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 421494 478102
rect 420874 477978 421494 478046
rect 420874 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 421494 477978
rect 420874 460350 421494 477922
rect 420874 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 421494 460350
rect 420874 460226 421494 460294
rect 420874 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 421494 460226
rect 420874 460102 421494 460170
rect 420874 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 421494 460102
rect 420874 459978 421494 460046
rect 420874 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 421494 459978
rect 420874 442350 421494 459922
rect 420874 442294 420970 442350
rect 421026 442294 421094 442350
rect 421150 442294 421218 442350
rect 421274 442294 421342 442350
rect 421398 442294 421494 442350
rect 420874 442226 421494 442294
rect 420874 442170 420970 442226
rect 421026 442170 421094 442226
rect 421150 442170 421218 442226
rect 421274 442170 421342 442226
rect 421398 442170 421494 442226
rect 420874 442102 421494 442170
rect 420874 442046 420970 442102
rect 421026 442046 421094 442102
rect 421150 442046 421218 442102
rect 421274 442046 421342 442102
rect 421398 442046 421494 442102
rect 420874 441978 421494 442046
rect 420874 441922 420970 441978
rect 421026 441922 421094 441978
rect 421150 441922 421218 441978
rect 421274 441922 421342 441978
rect 421398 441922 421494 441978
rect 402874 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 403494 424350
rect 402874 424226 403494 424294
rect 402874 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 403494 424226
rect 402874 424102 403494 424170
rect 402874 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 403494 424102
rect 402874 423978 403494 424046
rect 402874 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 403494 423978
rect 399154 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 399774 418350
rect 399154 418226 399774 418294
rect 399154 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 399774 418226
rect 399154 418102 399774 418170
rect 399154 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 399774 418102
rect 399154 417978 399774 418046
rect 399154 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 399774 417978
rect 384874 406294 384970 406350
rect 385026 406294 385094 406350
rect 385150 406294 385218 406350
rect 385274 406294 385342 406350
rect 385398 406294 385494 406350
rect 384874 406226 385494 406294
rect 384874 406170 384970 406226
rect 385026 406170 385094 406226
rect 385150 406170 385218 406226
rect 385274 406170 385342 406226
rect 385398 406170 385494 406226
rect 384874 406102 385494 406170
rect 384874 406046 384970 406102
rect 385026 406046 385094 406102
rect 385150 406046 385218 406102
rect 385274 406046 385342 406102
rect 385398 406046 385494 406102
rect 384874 405978 385494 406046
rect 384874 405922 384970 405978
rect 385026 405922 385094 405978
rect 385150 405922 385218 405978
rect 385274 405922 385342 405978
rect 385398 405922 385494 405978
rect 384874 388350 385494 405922
rect 387008 406350 387328 406384
rect 387008 406294 387078 406350
rect 387134 406294 387202 406350
rect 387258 406294 387328 406350
rect 387008 406226 387328 406294
rect 387008 406170 387078 406226
rect 387134 406170 387202 406226
rect 387258 406170 387328 406226
rect 387008 406102 387328 406170
rect 387008 406046 387078 406102
rect 387134 406046 387202 406102
rect 387258 406046 387328 406102
rect 387008 405978 387328 406046
rect 387008 405922 387078 405978
rect 387134 405922 387202 405978
rect 387258 405922 387328 405978
rect 387008 405888 387328 405922
rect 399154 400350 399774 417922
rect 402368 418350 402688 418384
rect 402368 418294 402438 418350
rect 402494 418294 402562 418350
rect 402618 418294 402688 418350
rect 402368 418226 402688 418294
rect 402368 418170 402438 418226
rect 402494 418170 402562 418226
rect 402618 418170 402688 418226
rect 402368 418102 402688 418170
rect 402368 418046 402438 418102
rect 402494 418046 402562 418102
rect 402618 418046 402688 418102
rect 402368 417978 402688 418046
rect 402368 417922 402438 417978
rect 402494 417922 402562 417978
rect 402618 417922 402688 417978
rect 402368 417888 402688 417922
rect 402874 406350 403494 423922
rect 417728 424350 418048 424384
rect 417728 424294 417798 424350
rect 417854 424294 417922 424350
rect 417978 424294 418048 424350
rect 417728 424226 418048 424294
rect 417728 424170 417798 424226
rect 417854 424170 417922 424226
rect 417978 424170 418048 424226
rect 417728 424102 418048 424170
rect 417728 424046 417798 424102
rect 417854 424046 417922 424102
rect 417978 424046 418048 424102
rect 417728 423978 418048 424046
rect 417728 423922 417798 423978
rect 417854 423922 417922 423978
rect 417978 423922 418048 423978
rect 417728 423888 418048 423922
rect 420874 424350 421494 441922
rect 435154 597212 435774 598268
rect 435154 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 435774 597212
rect 435154 597088 435774 597156
rect 435154 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 435774 597088
rect 435154 596964 435774 597032
rect 435154 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 435774 596964
rect 435154 596840 435774 596908
rect 435154 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 435774 596840
rect 435154 580350 435774 596784
rect 435154 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 435774 580350
rect 435154 580226 435774 580294
rect 435154 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 435774 580226
rect 435154 580102 435774 580170
rect 435154 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 435774 580102
rect 435154 579978 435774 580046
rect 435154 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 435774 579978
rect 435154 562350 435774 579922
rect 435154 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 435774 562350
rect 435154 562226 435774 562294
rect 435154 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 435774 562226
rect 435154 562102 435774 562170
rect 435154 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 435774 562102
rect 435154 561978 435774 562046
rect 435154 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 435774 561978
rect 435154 544350 435774 561922
rect 435154 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 435774 544350
rect 435154 544226 435774 544294
rect 435154 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 435774 544226
rect 435154 544102 435774 544170
rect 435154 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 435774 544102
rect 435154 543978 435774 544046
rect 435154 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 435774 543978
rect 435154 526350 435774 543922
rect 435154 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 435774 526350
rect 435154 526226 435774 526294
rect 435154 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 435774 526226
rect 435154 526102 435774 526170
rect 435154 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 435774 526102
rect 435154 525978 435774 526046
rect 435154 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 435774 525978
rect 435154 508350 435774 525922
rect 435154 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 435774 508350
rect 435154 508226 435774 508294
rect 435154 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 435774 508226
rect 435154 508102 435774 508170
rect 435154 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 435774 508102
rect 435154 507978 435774 508046
rect 435154 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 435774 507978
rect 435154 490350 435774 507922
rect 435154 490294 435250 490350
rect 435306 490294 435374 490350
rect 435430 490294 435498 490350
rect 435554 490294 435622 490350
rect 435678 490294 435774 490350
rect 435154 490226 435774 490294
rect 435154 490170 435250 490226
rect 435306 490170 435374 490226
rect 435430 490170 435498 490226
rect 435554 490170 435622 490226
rect 435678 490170 435774 490226
rect 435154 490102 435774 490170
rect 435154 490046 435250 490102
rect 435306 490046 435374 490102
rect 435430 490046 435498 490102
rect 435554 490046 435622 490102
rect 435678 490046 435774 490102
rect 435154 489978 435774 490046
rect 435154 489922 435250 489978
rect 435306 489922 435374 489978
rect 435430 489922 435498 489978
rect 435554 489922 435622 489978
rect 435678 489922 435774 489978
rect 435154 472350 435774 489922
rect 435154 472294 435250 472350
rect 435306 472294 435374 472350
rect 435430 472294 435498 472350
rect 435554 472294 435622 472350
rect 435678 472294 435774 472350
rect 435154 472226 435774 472294
rect 435154 472170 435250 472226
rect 435306 472170 435374 472226
rect 435430 472170 435498 472226
rect 435554 472170 435622 472226
rect 435678 472170 435774 472226
rect 435154 472102 435774 472170
rect 435154 472046 435250 472102
rect 435306 472046 435374 472102
rect 435430 472046 435498 472102
rect 435554 472046 435622 472102
rect 435678 472046 435774 472102
rect 435154 471978 435774 472046
rect 435154 471922 435250 471978
rect 435306 471922 435374 471978
rect 435430 471922 435498 471978
rect 435554 471922 435622 471978
rect 435678 471922 435774 471978
rect 435154 454350 435774 471922
rect 435154 454294 435250 454350
rect 435306 454294 435374 454350
rect 435430 454294 435498 454350
rect 435554 454294 435622 454350
rect 435678 454294 435774 454350
rect 435154 454226 435774 454294
rect 435154 454170 435250 454226
rect 435306 454170 435374 454226
rect 435430 454170 435498 454226
rect 435554 454170 435622 454226
rect 435678 454170 435774 454226
rect 435154 454102 435774 454170
rect 435154 454046 435250 454102
rect 435306 454046 435374 454102
rect 435430 454046 435498 454102
rect 435554 454046 435622 454102
rect 435678 454046 435774 454102
rect 435154 453978 435774 454046
rect 435154 453922 435250 453978
rect 435306 453922 435374 453978
rect 435430 453922 435498 453978
rect 435554 453922 435622 453978
rect 435678 453922 435774 453978
rect 433468 439348 433524 439358
rect 433468 438564 433524 439292
rect 433468 438498 433524 438508
rect 433088 436317 433408 436380
rect 433088 436261 433158 436317
rect 433214 436261 433282 436317
rect 433338 436261 433408 436317
rect 433088 436193 433408 436261
rect 433088 436137 433158 436193
rect 433214 436137 433282 436193
rect 433338 436137 433408 436193
rect 433088 436069 433408 436137
rect 433088 436013 433158 436069
rect 433214 436013 433282 436069
rect 433338 436013 433408 436069
rect 433088 435945 433408 436013
rect 433088 435889 433158 435945
rect 433214 435889 433282 435945
rect 433338 435889 433408 435945
rect 433088 435826 433408 435889
rect 435154 436350 435774 453922
rect 435154 436294 435250 436350
rect 435306 436294 435374 436350
rect 435430 436294 435498 436350
rect 435554 436294 435622 436350
rect 435678 436294 435774 436350
rect 435154 436226 435774 436294
rect 435154 436170 435250 436226
rect 435306 436170 435374 436226
rect 435430 436170 435498 436226
rect 435554 436170 435622 436226
rect 435678 436170 435774 436226
rect 435154 436102 435774 436170
rect 435154 436046 435250 436102
rect 435306 436046 435374 436102
rect 435430 436046 435498 436102
rect 435554 436046 435622 436102
rect 435678 436046 435774 436102
rect 435154 435978 435774 436046
rect 435154 435922 435250 435978
rect 435306 435922 435374 435978
rect 435430 435922 435498 435978
rect 435554 435922 435622 435978
rect 435678 435922 435774 435978
rect 420874 424294 420970 424350
rect 421026 424294 421094 424350
rect 421150 424294 421218 424350
rect 421274 424294 421342 424350
rect 421398 424294 421494 424350
rect 420874 424226 421494 424294
rect 420874 424170 420970 424226
rect 421026 424170 421094 424226
rect 421150 424170 421218 424226
rect 421274 424170 421342 424226
rect 421398 424170 421494 424226
rect 420874 424102 421494 424170
rect 420874 424046 420970 424102
rect 421026 424046 421094 424102
rect 421150 424046 421218 424102
rect 421274 424046 421342 424102
rect 421398 424046 421494 424102
rect 420874 423978 421494 424046
rect 420874 423922 420970 423978
rect 421026 423922 421094 423978
rect 421150 423922 421218 423978
rect 421274 423922 421342 423978
rect 421398 423922 421494 423978
rect 402874 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 403494 406350
rect 402874 406226 403494 406294
rect 402874 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 403494 406226
rect 402874 406102 403494 406170
rect 402874 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 403494 406102
rect 402874 405978 403494 406046
rect 402874 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 403494 405978
rect 399154 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 399774 400350
rect 399154 400226 399774 400294
rect 399154 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 399774 400226
rect 399154 400102 399774 400170
rect 399154 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 399774 400102
rect 399154 399978 399774 400046
rect 399154 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 399774 399978
rect 384874 388294 384970 388350
rect 385026 388294 385094 388350
rect 385150 388294 385218 388350
rect 385274 388294 385342 388350
rect 385398 388294 385494 388350
rect 384874 388226 385494 388294
rect 384874 388170 384970 388226
rect 385026 388170 385094 388226
rect 385150 388170 385218 388226
rect 385274 388170 385342 388226
rect 385398 388170 385494 388226
rect 384874 388102 385494 388170
rect 384874 388046 384970 388102
rect 385026 388046 385094 388102
rect 385150 388046 385218 388102
rect 385274 388046 385342 388102
rect 385398 388046 385494 388102
rect 384874 387978 385494 388046
rect 384874 387922 384970 387978
rect 385026 387922 385094 387978
rect 385150 387922 385218 387978
rect 385274 387922 385342 387978
rect 385398 387922 385494 387978
rect 384874 370350 385494 387922
rect 387008 388350 387328 388384
rect 387008 388294 387078 388350
rect 387134 388294 387202 388350
rect 387258 388294 387328 388350
rect 387008 388226 387328 388294
rect 387008 388170 387078 388226
rect 387134 388170 387202 388226
rect 387258 388170 387328 388226
rect 387008 388102 387328 388170
rect 387008 388046 387078 388102
rect 387134 388046 387202 388102
rect 387258 388046 387328 388102
rect 387008 387978 387328 388046
rect 387008 387922 387078 387978
rect 387134 387922 387202 387978
rect 387258 387922 387328 387978
rect 387008 387888 387328 387922
rect 399154 382350 399774 399922
rect 402368 400350 402688 400384
rect 402368 400294 402438 400350
rect 402494 400294 402562 400350
rect 402618 400294 402688 400350
rect 402368 400226 402688 400294
rect 402368 400170 402438 400226
rect 402494 400170 402562 400226
rect 402618 400170 402688 400226
rect 402368 400102 402688 400170
rect 402368 400046 402438 400102
rect 402494 400046 402562 400102
rect 402618 400046 402688 400102
rect 402368 399978 402688 400046
rect 402368 399922 402438 399978
rect 402494 399922 402562 399978
rect 402618 399922 402688 399978
rect 402368 399888 402688 399922
rect 402874 388350 403494 405922
rect 417728 406350 418048 406384
rect 417728 406294 417798 406350
rect 417854 406294 417922 406350
rect 417978 406294 418048 406350
rect 417728 406226 418048 406294
rect 417728 406170 417798 406226
rect 417854 406170 417922 406226
rect 417978 406170 418048 406226
rect 417728 406102 418048 406170
rect 417728 406046 417798 406102
rect 417854 406046 417922 406102
rect 417978 406046 418048 406102
rect 417728 405978 418048 406046
rect 417728 405922 417798 405978
rect 417854 405922 417922 405978
rect 417978 405922 418048 405978
rect 417728 405888 418048 405922
rect 420874 406350 421494 423922
rect 433088 418350 433408 418384
rect 433088 418294 433158 418350
rect 433214 418294 433282 418350
rect 433338 418294 433408 418350
rect 433088 418226 433408 418294
rect 433088 418170 433158 418226
rect 433214 418170 433282 418226
rect 433338 418170 433408 418226
rect 433088 418102 433408 418170
rect 433088 418046 433158 418102
rect 433214 418046 433282 418102
rect 433338 418046 433408 418102
rect 433088 417978 433408 418046
rect 433088 417922 433158 417978
rect 433214 417922 433282 417978
rect 433338 417922 433408 417978
rect 433088 417888 433408 417922
rect 435154 418350 435774 435922
rect 435154 418294 435250 418350
rect 435306 418294 435374 418350
rect 435430 418294 435498 418350
rect 435554 418294 435622 418350
rect 435678 418294 435774 418350
rect 435154 418226 435774 418294
rect 435154 418170 435250 418226
rect 435306 418170 435374 418226
rect 435430 418170 435498 418226
rect 435554 418170 435622 418226
rect 435678 418170 435774 418226
rect 435154 418102 435774 418170
rect 435154 418046 435250 418102
rect 435306 418046 435374 418102
rect 435430 418046 435498 418102
rect 435554 418046 435622 418102
rect 435678 418046 435774 418102
rect 435154 417978 435774 418046
rect 435154 417922 435250 417978
rect 435306 417922 435374 417978
rect 435430 417922 435498 417978
rect 435554 417922 435622 417978
rect 435678 417922 435774 417978
rect 420874 406294 420970 406350
rect 421026 406294 421094 406350
rect 421150 406294 421218 406350
rect 421274 406294 421342 406350
rect 421398 406294 421494 406350
rect 420874 406226 421494 406294
rect 420874 406170 420970 406226
rect 421026 406170 421094 406226
rect 421150 406170 421218 406226
rect 421274 406170 421342 406226
rect 421398 406170 421494 406226
rect 420874 406102 421494 406170
rect 420874 406046 420970 406102
rect 421026 406046 421094 406102
rect 421150 406046 421218 406102
rect 421274 406046 421342 406102
rect 421398 406046 421494 406102
rect 420874 405978 421494 406046
rect 420874 405922 420970 405978
rect 421026 405922 421094 405978
rect 421150 405922 421218 405978
rect 421274 405922 421342 405978
rect 421398 405922 421494 405978
rect 402874 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 403494 388350
rect 402874 388226 403494 388294
rect 402874 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 403494 388226
rect 402874 388102 403494 388170
rect 402874 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 403494 388102
rect 402874 387978 403494 388046
rect 402874 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 403494 387978
rect 399154 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 399774 382350
rect 399154 382226 399774 382294
rect 399154 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 399774 382226
rect 399154 382102 399774 382170
rect 399154 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 399774 382102
rect 399154 381978 399774 382046
rect 399154 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 399774 381978
rect 384874 370294 384970 370350
rect 385026 370294 385094 370350
rect 385150 370294 385218 370350
rect 385274 370294 385342 370350
rect 385398 370294 385494 370350
rect 384874 370226 385494 370294
rect 384874 370170 384970 370226
rect 385026 370170 385094 370226
rect 385150 370170 385218 370226
rect 385274 370170 385342 370226
rect 385398 370170 385494 370226
rect 384874 370102 385494 370170
rect 384874 370046 384970 370102
rect 385026 370046 385094 370102
rect 385150 370046 385218 370102
rect 385274 370046 385342 370102
rect 385398 370046 385494 370102
rect 384874 369978 385494 370046
rect 384874 369922 384970 369978
rect 385026 369922 385094 369978
rect 385150 369922 385218 369978
rect 385274 369922 385342 369978
rect 385398 369922 385494 369978
rect 384874 352350 385494 369922
rect 387008 370350 387328 370384
rect 387008 370294 387078 370350
rect 387134 370294 387202 370350
rect 387258 370294 387328 370350
rect 387008 370226 387328 370294
rect 387008 370170 387078 370226
rect 387134 370170 387202 370226
rect 387258 370170 387328 370226
rect 387008 370102 387328 370170
rect 387008 370046 387078 370102
rect 387134 370046 387202 370102
rect 387258 370046 387328 370102
rect 387008 369978 387328 370046
rect 387008 369922 387078 369978
rect 387134 369922 387202 369978
rect 387258 369922 387328 369978
rect 387008 369888 387328 369922
rect 399154 364350 399774 381922
rect 402368 382350 402688 382384
rect 402368 382294 402438 382350
rect 402494 382294 402562 382350
rect 402618 382294 402688 382350
rect 402368 382226 402688 382294
rect 402368 382170 402438 382226
rect 402494 382170 402562 382226
rect 402618 382170 402688 382226
rect 402368 382102 402688 382170
rect 402368 382046 402438 382102
rect 402494 382046 402562 382102
rect 402618 382046 402688 382102
rect 402368 381978 402688 382046
rect 402368 381922 402438 381978
rect 402494 381922 402562 381978
rect 402618 381922 402688 381978
rect 402368 381888 402688 381922
rect 402874 370350 403494 387922
rect 417728 388350 418048 388384
rect 417728 388294 417798 388350
rect 417854 388294 417922 388350
rect 417978 388294 418048 388350
rect 417728 388226 418048 388294
rect 417728 388170 417798 388226
rect 417854 388170 417922 388226
rect 417978 388170 418048 388226
rect 417728 388102 418048 388170
rect 417728 388046 417798 388102
rect 417854 388046 417922 388102
rect 417978 388046 418048 388102
rect 417728 387978 418048 388046
rect 417728 387922 417798 387978
rect 417854 387922 417922 387978
rect 417978 387922 418048 387978
rect 417728 387888 418048 387922
rect 420874 388350 421494 405922
rect 433088 400350 433408 400384
rect 433088 400294 433158 400350
rect 433214 400294 433282 400350
rect 433338 400294 433408 400350
rect 433088 400226 433408 400294
rect 433088 400170 433158 400226
rect 433214 400170 433282 400226
rect 433338 400170 433408 400226
rect 433088 400102 433408 400170
rect 433088 400046 433158 400102
rect 433214 400046 433282 400102
rect 433338 400046 433408 400102
rect 433088 399978 433408 400046
rect 433088 399922 433158 399978
rect 433214 399922 433282 399978
rect 433338 399922 433408 399978
rect 433088 399888 433408 399922
rect 435154 400350 435774 417922
rect 435154 400294 435250 400350
rect 435306 400294 435374 400350
rect 435430 400294 435498 400350
rect 435554 400294 435622 400350
rect 435678 400294 435774 400350
rect 435154 400226 435774 400294
rect 435154 400170 435250 400226
rect 435306 400170 435374 400226
rect 435430 400170 435498 400226
rect 435554 400170 435622 400226
rect 435678 400170 435774 400226
rect 435154 400102 435774 400170
rect 435154 400046 435250 400102
rect 435306 400046 435374 400102
rect 435430 400046 435498 400102
rect 435554 400046 435622 400102
rect 435678 400046 435774 400102
rect 435154 399978 435774 400046
rect 435154 399922 435250 399978
rect 435306 399922 435374 399978
rect 435430 399922 435498 399978
rect 435554 399922 435622 399978
rect 435678 399922 435774 399978
rect 420874 388294 420970 388350
rect 421026 388294 421094 388350
rect 421150 388294 421218 388350
rect 421274 388294 421342 388350
rect 421398 388294 421494 388350
rect 420874 388226 421494 388294
rect 420874 388170 420970 388226
rect 421026 388170 421094 388226
rect 421150 388170 421218 388226
rect 421274 388170 421342 388226
rect 421398 388170 421494 388226
rect 420874 388102 421494 388170
rect 420874 388046 420970 388102
rect 421026 388046 421094 388102
rect 421150 388046 421218 388102
rect 421274 388046 421342 388102
rect 421398 388046 421494 388102
rect 420874 387978 421494 388046
rect 420874 387922 420970 387978
rect 421026 387922 421094 387978
rect 421150 387922 421218 387978
rect 421274 387922 421342 387978
rect 421398 387922 421494 387978
rect 402874 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 403494 370350
rect 402874 370226 403494 370294
rect 402874 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 403494 370226
rect 402874 370102 403494 370170
rect 402874 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 403494 370102
rect 402874 369978 403494 370046
rect 402874 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 403494 369978
rect 399154 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 399774 364350
rect 399154 364226 399774 364294
rect 399154 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 399774 364226
rect 399154 364102 399774 364170
rect 399154 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 399774 364102
rect 399154 363978 399774 364046
rect 399154 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 399774 363978
rect 384874 352294 384970 352350
rect 385026 352294 385094 352350
rect 385150 352294 385218 352350
rect 385274 352294 385342 352350
rect 385398 352294 385494 352350
rect 384874 352226 385494 352294
rect 384874 352170 384970 352226
rect 385026 352170 385094 352226
rect 385150 352170 385218 352226
rect 385274 352170 385342 352226
rect 385398 352170 385494 352226
rect 384874 352102 385494 352170
rect 384874 352046 384970 352102
rect 385026 352046 385094 352102
rect 385150 352046 385218 352102
rect 385274 352046 385342 352102
rect 385398 352046 385494 352102
rect 384874 351978 385494 352046
rect 384874 351922 384970 351978
rect 385026 351922 385094 351978
rect 385150 351922 385218 351978
rect 385274 351922 385342 351978
rect 385398 351922 385494 351978
rect 384874 334350 385494 351922
rect 387008 352350 387328 352384
rect 387008 352294 387078 352350
rect 387134 352294 387202 352350
rect 387258 352294 387328 352350
rect 387008 352226 387328 352294
rect 387008 352170 387078 352226
rect 387134 352170 387202 352226
rect 387258 352170 387328 352226
rect 387008 352102 387328 352170
rect 387008 352046 387078 352102
rect 387134 352046 387202 352102
rect 387258 352046 387328 352102
rect 387008 351978 387328 352046
rect 387008 351922 387078 351978
rect 387134 351922 387202 351978
rect 387258 351922 387328 351978
rect 387008 351888 387328 351922
rect 399154 346350 399774 363922
rect 402368 364350 402688 364384
rect 402368 364294 402438 364350
rect 402494 364294 402562 364350
rect 402618 364294 402688 364350
rect 402368 364226 402688 364294
rect 402368 364170 402438 364226
rect 402494 364170 402562 364226
rect 402618 364170 402688 364226
rect 402368 364102 402688 364170
rect 402368 364046 402438 364102
rect 402494 364046 402562 364102
rect 402618 364046 402688 364102
rect 402368 363978 402688 364046
rect 402368 363922 402438 363978
rect 402494 363922 402562 363978
rect 402618 363922 402688 363978
rect 402368 363888 402688 363922
rect 402874 352350 403494 369922
rect 417728 370350 418048 370384
rect 417728 370294 417798 370350
rect 417854 370294 417922 370350
rect 417978 370294 418048 370350
rect 417728 370226 418048 370294
rect 417728 370170 417798 370226
rect 417854 370170 417922 370226
rect 417978 370170 418048 370226
rect 417728 370102 418048 370170
rect 417728 370046 417798 370102
rect 417854 370046 417922 370102
rect 417978 370046 418048 370102
rect 417728 369978 418048 370046
rect 417728 369922 417798 369978
rect 417854 369922 417922 369978
rect 417978 369922 418048 369978
rect 417728 369888 418048 369922
rect 420874 370350 421494 387922
rect 433088 382350 433408 382384
rect 433088 382294 433158 382350
rect 433214 382294 433282 382350
rect 433338 382294 433408 382350
rect 433088 382226 433408 382294
rect 433088 382170 433158 382226
rect 433214 382170 433282 382226
rect 433338 382170 433408 382226
rect 433088 382102 433408 382170
rect 433088 382046 433158 382102
rect 433214 382046 433282 382102
rect 433338 382046 433408 382102
rect 433088 381978 433408 382046
rect 433088 381922 433158 381978
rect 433214 381922 433282 381978
rect 433338 381922 433408 381978
rect 433088 381888 433408 381922
rect 435154 382350 435774 399922
rect 435154 382294 435250 382350
rect 435306 382294 435374 382350
rect 435430 382294 435498 382350
rect 435554 382294 435622 382350
rect 435678 382294 435774 382350
rect 435154 382226 435774 382294
rect 435154 382170 435250 382226
rect 435306 382170 435374 382226
rect 435430 382170 435498 382226
rect 435554 382170 435622 382226
rect 435678 382170 435774 382226
rect 435154 382102 435774 382170
rect 435154 382046 435250 382102
rect 435306 382046 435374 382102
rect 435430 382046 435498 382102
rect 435554 382046 435622 382102
rect 435678 382046 435774 382102
rect 435154 381978 435774 382046
rect 435154 381922 435250 381978
rect 435306 381922 435374 381978
rect 435430 381922 435498 381978
rect 435554 381922 435622 381978
rect 435678 381922 435774 381978
rect 420874 370294 420970 370350
rect 421026 370294 421094 370350
rect 421150 370294 421218 370350
rect 421274 370294 421342 370350
rect 421398 370294 421494 370350
rect 420874 370226 421494 370294
rect 420874 370170 420970 370226
rect 421026 370170 421094 370226
rect 421150 370170 421218 370226
rect 421274 370170 421342 370226
rect 421398 370170 421494 370226
rect 420874 370102 421494 370170
rect 420874 370046 420970 370102
rect 421026 370046 421094 370102
rect 421150 370046 421218 370102
rect 421274 370046 421342 370102
rect 421398 370046 421494 370102
rect 420874 369978 421494 370046
rect 420874 369922 420970 369978
rect 421026 369922 421094 369978
rect 421150 369922 421218 369978
rect 421274 369922 421342 369978
rect 421398 369922 421494 369978
rect 402874 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 403494 352350
rect 402874 352226 403494 352294
rect 402874 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 403494 352226
rect 402874 352102 403494 352170
rect 402874 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 403494 352102
rect 402874 351978 403494 352046
rect 402874 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 403494 351978
rect 399154 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 399774 346350
rect 399154 346226 399774 346294
rect 399154 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 399774 346226
rect 399154 346102 399774 346170
rect 399154 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 399774 346102
rect 399154 345978 399774 346046
rect 399154 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 399774 345978
rect 384874 334294 384970 334350
rect 385026 334294 385094 334350
rect 385150 334294 385218 334350
rect 385274 334294 385342 334350
rect 385398 334294 385494 334350
rect 384874 334226 385494 334294
rect 384874 334170 384970 334226
rect 385026 334170 385094 334226
rect 385150 334170 385218 334226
rect 385274 334170 385342 334226
rect 385398 334170 385494 334226
rect 384874 334102 385494 334170
rect 384874 334046 384970 334102
rect 385026 334046 385094 334102
rect 385150 334046 385218 334102
rect 385274 334046 385342 334102
rect 385398 334046 385494 334102
rect 384874 333978 385494 334046
rect 384874 333922 384970 333978
rect 385026 333922 385094 333978
rect 385150 333922 385218 333978
rect 385274 333922 385342 333978
rect 385398 333922 385494 333978
rect 384874 316350 385494 333922
rect 387008 334350 387328 334384
rect 387008 334294 387078 334350
rect 387134 334294 387202 334350
rect 387258 334294 387328 334350
rect 387008 334226 387328 334294
rect 387008 334170 387078 334226
rect 387134 334170 387202 334226
rect 387258 334170 387328 334226
rect 387008 334102 387328 334170
rect 387008 334046 387078 334102
rect 387134 334046 387202 334102
rect 387258 334046 387328 334102
rect 387008 333978 387328 334046
rect 387008 333922 387078 333978
rect 387134 333922 387202 333978
rect 387258 333922 387328 333978
rect 387008 333888 387328 333922
rect 399154 328350 399774 345922
rect 402368 346350 402688 346384
rect 402368 346294 402438 346350
rect 402494 346294 402562 346350
rect 402618 346294 402688 346350
rect 402368 346226 402688 346294
rect 402368 346170 402438 346226
rect 402494 346170 402562 346226
rect 402618 346170 402688 346226
rect 402368 346102 402688 346170
rect 402368 346046 402438 346102
rect 402494 346046 402562 346102
rect 402618 346046 402688 346102
rect 402368 345978 402688 346046
rect 402368 345922 402438 345978
rect 402494 345922 402562 345978
rect 402618 345922 402688 345978
rect 402368 345888 402688 345922
rect 402874 334350 403494 351922
rect 417728 352350 418048 352384
rect 417728 352294 417798 352350
rect 417854 352294 417922 352350
rect 417978 352294 418048 352350
rect 417728 352226 418048 352294
rect 417728 352170 417798 352226
rect 417854 352170 417922 352226
rect 417978 352170 418048 352226
rect 417728 352102 418048 352170
rect 417728 352046 417798 352102
rect 417854 352046 417922 352102
rect 417978 352046 418048 352102
rect 417728 351978 418048 352046
rect 417728 351922 417798 351978
rect 417854 351922 417922 351978
rect 417978 351922 418048 351978
rect 417728 351888 418048 351922
rect 420874 352350 421494 369922
rect 433088 364350 433408 364384
rect 433088 364294 433158 364350
rect 433214 364294 433282 364350
rect 433338 364294 433408 364350
rect 433088 364226 433408 364294
rect 433088 364170 433158 364226
rect 433214 364170 433282 364226
rect 433338 364170 433408 364226
rect 433088 364102 433408 364170
rect 433088 364046 433158 364102
rect 433214 364046 433282 364102
rect 433338 364046 433408 364102
rect 433088 363978 433408 364046
rect 433088 363922 433158 363978
rect 433214 363922 433282 363978
rect 433338 363922 433408 363978
rect 433088 363888 433408 363922
rect 435154 364350 435774 381922
rect 435154 364294 435250 364350
rect 435306 364294 435374 364350
rect 435430 364294 435498 364350
rect 435554 364294 435622 364350
rect 435678 364294 435774 364350
rect 435154 364226 435774 364294
rect 435154 364170 435250 364226
rect 435306 364170 435374 364226
rect 435430 364170 435498 364226
rect 435554 364170 435622 364226
rect 435678 364170 435774 364226
rect 435154 364102 435774 364170
rect 435154 364046 435250 364102
rect 435306 364046 435374 364102
rect 435430 364046 435498 364102
rect 435554 364046 435622 364102
rect 435678 364046 435774 364102
rect 435154 363978 435774 364046
rect 435154 363922 435250 363978
rect 435306 363922 435374 363978
rect 435430 363922 435498 363978
rect 435554 363922 435622 363978
rect 435678 363922 435774 363978
rect 420874 352294 420970 352350
rect 421026 352294 421094 352350
rect 421150 352294 421218 352350
rect 421274 352294 421342 352350
rect 421398 352294 421494 352350
rect 420874 352226 421494 352294
rect 420874 352170 420970 352226
rect 421026 352170 421094 352226
rect 421150 352170 421218 352226
rect 421274 352170 421342 352226
rect 421398 352170 421494 352226
rect 420874 352102 421494 352170
rect 420874 352046 420970 352102
rect 421026 352046 421094 352102
rect 421150 352046 421218 352102
rect 421274 352046 421342 352102
rect 421398 352046 421494 352102
rect 420874 351978 421494 352046
rect 420874 351922 420970 351978
rect 421026 351922 421094 351978
rect 421150 351922 421218 351978
rect 421274 351922 421342 351978
rect 421398 351922 421494 351978
rect 402874 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 403494 334350
rect 402874 334226 403494 334294
rect 402874 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 403494 334226
rect 402874 334102 403494 334170
rect 402874 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 403494 334102
rect 402874 333978 403494 334046
rect 402874 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 403494 333978
rect 399154 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 399774 328350
rect 399154 328226 399774 328294
rect 399154 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 399774 328226
rect 399154 328102 399774 328170
rect 399154 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 399774 328102
rect 399154 327978 399774 328046
rect 399154 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 399774 327978
rect 384874 316294 384970 316350
rect 385026 316294 385094 316350
rect 385150 316294 385218 316350
rect 385274 316294 385342 316350
rect 385398 316294 385494 316350
rect 384874 316226 385494 316294
rect 384874 316170 384970 316226
rect 385026 316170 385094 316226
rect 385150 316170 385218 316226
rect 385274 316170 385342 316226
rect 385398 316170 385494 316226
rect 384874 316102 385494 316170
rect 384874 316046 384970 316102
rect 385026 316046 385094 316102
rect 385150 316046 385218 316102
rect 385274 316046 385342 316102
rect 385398 316046 385494 316102
rect 384874 315978 385494 316046
rect 384874 315922 384970 315978
rect 385026 315922 385094 315978
rect 385150 315922 385218 315978
rect 385274 315922 385342 315978
rect 385398 315922 385494 315978
rect 384874 298350 385494 315922
rect 387008 316350 387328 316384
rect 387008 316294 387078 316350
rect 387134 316294 387202 316350
rect 387258 316294 387328 316350
rect 387008 316226 387328 316294
rect 387008 316170 387078 316226
rect 387134 316170 387202 316226
rect 387258 316170 387328 316226
rect 387008 316102 387328 316170
rect 387008 316046 387078 316102
rect 387134 316046 387202 316102
rect 387258 316046 387328 316102
rect 387008 315978 387328 316046
rect 387008 315922 387078 315978
rect 387134 315922 387202 315978
rect 387258 315922 387328 315978
rect 387008 315888 387328 315922
rect 399154 310350 399774 327922
rect 402368 328350 402688 328384
rect 402368 328294 402438 328350
rect 402494 328294 402562 328350
rect 402618 328294 402688 328350
rect 402368 328226 402688 328294
rect 402368 328170 402438 328226
rect 402494 328170 402562 328226
rect 402618 328170 402688 328226
rect 402368 328102 402688 328170
rect 402368 328046 402438 328102
rect 402494 328046 402562 328102
rect 402618 328046 402688 328102
rect 402368 327978 402688 328046
rect 402368 327922 402438 327978
rect 402494 327922 402562 327978
rect 402618 327922 402688 327978
rect 402368 327888 402688 327922
rect 402874 316350 403494 333922
rect 417728 334350 418048 334384
rect 417728 334294 417798 334350
rect 417854 334294 417922 334350
rect 417978 334294 418048 334350
rect 417728 334226 418048 334294
rect 417728 334170 417798 334226
rect 417854 334170 417922 334226
rect 417978 334170 418048 334226
rect 417728 334102 418048 334170
rect 417728 334046 417798 334102
rect 417854 334046 417922 334102
rect 417978 334046 418048 334102
rect 417728 333978 418048 334046
rect 417728 333922 417798 333978
rect 417854 333922 417922 333978
rect 417978 333922 418048 333978
rect 417728 333888 418048 333922
rect 420874 334350 421494 351922
rect 433088 346350 433408 346384
rect 433088 346294 433158 346350
rect 433214 346294 433282 346350
rect 433338 346294 433408 346350
rect 433088 346226 433408 346294
rect 433088 346170 433158 346226
rect 433214 346170 433282 346226
rect 433338 346170 433408 346226
rect 433088 346102 433408 346170
rect 433088 346046 433158 346102
rect 433214 346046 433282 346102
rect 433338 346046 433408 346102
rect 433088 345978 433408 346046
rect 433088 345922 433158 345978
rect 433214 345922 433282 345978
rect 433338 345922 433408 345978
rect 433088 345888 433408 345922
rect 435154 346350 435774 363922
rect 435154 346294 435250 346350
rect 435306 346294 435374 346350
rect 435430 346294 435498 346350
rect 435554 346294 435622 346350
rect 435678 346294 435774 346350
rect 435154 346226 435774 346294
rect 435154 346170 435250 346226
rect 435306 346170 435374 346226
rect 435430 346170 435498 346226
rect 435554 346170 435622 346226
rect 435678 346170 435774 346226
rect 435154 346102 435774 346170
rect 435154 346046 435250 346102
rect 435306 346046 435374 346102
rect 435430 346046 435498 346102
rect 435554 346046 435622 346102
rect 435678 346046 435774 346102
rect 435154 345978 435774 346046
rect 435154 345922 435250 345978
rect 435306 345922 435374 345978
rect 435430 345922 435498 345978
rect 435554 345922 435622 345978
rect 435678 345922 435774 345978
rect 420874 334294 420970 334350
rect 421026 334294 421094 334350
rect 421150 334294 421218 334350
rect 421274 334294 421342 334350
rect 421398 334294 421494 334350
rect 420874 334226 421494 334294
rect 420874 334170 420970 334226
rect 421026 334170 421094 334226
rect 421150 334170 421218 334226
rect 421274 334170 421342 334226
rect 421398 334170 421494 334226
rect 420874 334102 421494 334170
rect 420874 334046 420970 334102
rect 421026 334046 421094 334102
rect 421150 334046 421218 334102
rect 421274 334046 421342 334102
rect 421398 334046 421494 334102
rect 420874 333978 421494 334046
rect 420874 333922 420970 333978
rect 421026 333922 421094 333978
rect 421150 333922 421218 333978
rect 421274 333922 421342 333978
rect 421398 333922 421494 333978
rect 402874 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 403494 316350
rect 402874 316226 403494 316294
rect 402874 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 403494 316226
rect 402874 316102 403494 316170
rect 402874 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 403494 316102
rect 402874 315978 403494 316046
rect 402874 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 403494 315978
rect 399154 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 399774 310350
rect 399154 310226 399774 310294
rect 399154 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 399774 310226
rect 399154 310102 399774 310170
rect 399154 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 399774 310102
rect 399154 309978 399774 310046
rect 399154 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 399774 309978
rect 384874 298294 384970 298350
rect 385026 298294 385094 298350
rect 385150 298294 385218 298350
rect 385274 298294 385342 298350
rect 385398 298294 385494 298350
rect 384874 298226 385494 298294
rect 384874 298170 384970 298226
rect 385026 298170 385094 298226
rect 385150 298170 385218 298226
rect 385274 298170 385342 298226
rect 385398 298170 385494 298226
rect 384874 298102 385494 298170
rect 384874 298046 384970 298102
rect 385026 298046 385094 298102
rect 385150 298046 385218 298102
rect 385274 298046 385342 298102
rect 385398 298046 385494 298102
rect 384874 297978 385494 298046
rect 384874 297922 384970 297978
rect 385026 297922 385094 297978
rect 385150 297922 385218 297978
rect 385274 297922 385342 297978
rect 385398 297922 385494 297978
rect 384874 280350 385494 297922
rect 387008 298350 387328 298384
rect 387008 298294 387078 298350
rect 387134 298294 387202 298350
rect 387258 298294 387328 298350
rect 387008 298226 387328 298294
rect 387008 298170 387078 298226
rect 387134 298170 387202 298226
rect 387258 298170 387328 298226
rect 387008 298102 387328 298170
rect 387008 298046 387078 298102
rect 387134 298046 387202 298102
rect 387258 298046 387328 298102
rect 387008 297978 387328 298046
rect 387008 297922 387078 297978
rect 387134 297922 387202 297978
rect 387258 297922 387328 297978
rect 387008 297888 387328 297922
rect 399154 292350 399774 309922
rect 402368 310350 402688 310384
rect 402368 310294 402438 310350
rect 402494 310294 402562 310350
rect 402618 310294 402688 310350
rect 402368 310226 402688 310294
rect 402368 310170 402438 310226
rect 402494 310170 402562 310226
rect 402618 310170 402688 310226
rect 402368 310102 402688 310170
rect 402368 310046 402438 310102
rect 402494 310046 402562 310102
rect 402618 310046 402688 310102
rect 402368 309978 402688 310046
rect 402368 309922 402438 309978
rect 402494 309922 402562 309978
rect 402618 309922 402688 309978
rect 402368 309888 402688 309922
rect 402874 298350 403494 315922
rect 417728 316350 418048 316384
rect 417728 316294 417798 316350
rect 417854 316294 417922 316350
rect 417978 316294 418048 316350
rect 417728 316226 418048 316294
rect 417728 316170 417798 316226
rect 417854 316170 417922 316226
rect 417978 316170 418048 316226
rect 417728 316102 418048 316170
rect 417728 316046 417798 316102
rect 417854 316046 417922 316102
rect 417978 316046 418048 316102
rect 417728 315978 418048 316046
rect 417728 315922 417798 315978
rect 417854 315922 417922 315978
rect 417978 315922 418048 315978
rect 417728 315888 418048 315922
rect 420874 316350 421494 333922
rect 433088 328350 433408 328384
rect 433088 328294 433158 328350
rect 433214 328294 433282 328350
rect 433338 328294 433408 328350
rect 433088 328226 433408 328294
rect 433088 328170 433158 328226
rect 433214 328170 433282 328226
rect 433338 328170 433408 328226
rect 433088 328102 433408 328170
rect 433088 328046 433158 328102
rect 433214 328046 433282 328102
rect 433338 328046 433408 328102
rect 433088 327978 433408 328046
rect 433088 327922 433158 327978
rect 433214 327922 433282 327978
rect 433338 327922 433408 327978
rect 433088 327888 433408 327922
rect 435154 328350 435774 345922
rect 435154 328294 435250 328350
rect 435306 328294 435374 328350
rect 435430 328294 435498 328350
rect 435554 328294 435622 328350
rect 435678 328294 435774 328350
rect 435154 328226 435774 328294
rect 435154 328170 435250 328226
rect 435306 328170 435374 328226
rect 435430 328170 435498 328226
rect 435554 328170 435622 328226
rect 435678 328170 435774 328226
rect 435154 328102 435774 328170
rect 435154 328046 435250 328102
rect 435306 328046 435374 328102
rect 435430 328046 435498 328102
rect 435554 328046 435622 328102
rect 435678 328046 435774 328102
rect 435154 327978 435774 328046
rect 435154 327922 435250 327978
rect 435306 327922 435374 327978
rect 435430 327922 435498 327978
rect 435554 327922 435622 327978
rect 435678 327922 435774 327978
rect 420874 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 421494 316350
rect 420874 316226 421494 316294
rect 420874 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 421494 316226
rect 420874 316102 421494 316170
rect 420874 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 421494 316102
rect 420874 315978 421494 316046
rect 420874 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 421494 315978
rect 402874 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 403494 298350
rect 402874 298226 403494 298294
rect 402874 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 403494 298226
rect 402874 298102 403494 298170
rect 402874 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 403494 298102
rect 402874 297978 403494 298046
rect 402874 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 403494 297978
rect 399154 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 399774 292350
rect 399154 292226 399774 292294
rect 399154 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 399774 292226
rect 399154 292102 399774 292170
rect 399154 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 399774 292102
rect 399154 291978 399774 292046
rect 399154 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 399774 291978
rect 384874 280294 384970 280350
rect 385026 280294 385094 280350
rect 385150 280294 385218 280350
rect 385274 280294 385342 280350
rect 385398 280294 385494 280350
rect 384874 280226 385494 280294
rect 384874 280170 384970 280226
rect 385026 280170 385094 280226
rect 385150 280170 385218 280226
rect 385274 280170 385342 280226
rect 385398 280170 385494 280226
rect 384874 280102 385494 280170
rect 384874 280046 384970 280102
rect 385026 280046 385094 280102
rect 385150 280046 385218 280102
rect 385274 280046 385342 280102
rect 385398 280046 385494 280102
rect 384874 279978 385494 280046
rect 384874 279922 384970 279978
rect 385026 279922 385094 279978
rect 385150 279922 385218 279978
rect 385274 279922 385342 279978
rect 385398 279922 385494 279978
rect 384874 262350 385494 279922
rect 387008 280350 387328 280384
rect 387008 280294 387078 280350
rect 387134 280294 387202 280350
rect 387258 280294 387328 280350
rect 387008 280226 387328 280294
rect 387008 280170 387078 280226
rect 387134 280170 387202 280226
rect 387258 280170 387328 280226
rect 387008 280102 387328 280170
rect 387008 280046 387078 280102
rect 387134 280046 387202 280102
rect 387258 280046 387328 280102
rect 387008 279978 387328 280046
rect 387008 279922 387078 279978
rect 387134 279922 387202 279978
rect 387258 279922 387328 279978
rect 387008 279888 387328 279922
rect 399154 274350 399774 291922
rect 402368 292350 402688 292384
rect 402368 292294 402438 292350
rect 402494 292294 402562 292350
rect 402618 292294 402688 292350
rect 402368 292226 402688 292294
rect 402368 292170 402438 292226
rect 402494 292170 402562 292226
rect 402618 292170 402688 292226
rect 402368 292102 402688 292170
rect 402368 292046 402438 292102
rect 402494 292046 402562 292102
rect 402618 292046 402688 292102
rect 402368 291978 402688 292046
rect 402368 291922 402438 291978
rect 402494 291922 402562 291978
rect 402618 291922 402688 291978
rect 402368 291888 402688 291922
rect 402874 280350 403494 297922
rect 417728 298350 418048 298384
rect 417728 298294 417798 298350
rect 417854 298294 417922 298350
rect 417978 298294 418048 298350
rect 417728 298226 418048 298294
rect 417728 298170 417798 298226
rect 417854 298170 417922 298226
rect 417978 298170 418048 298226
rect 417728 298102 418048 298170
rect 417728 298046 417798 298102
rect 417854 298046 417922 298102
rect 417978 298046 418048 298102
rect 417728 297978 418048 298046
rect 417728 297922 417798 297978
rect 417854 297922 417922 297978
rect 417978 297922 418048 297978
rect 417728 297888 418048 297922
rect 420874 298350 421494 315922
rect 433088 310350 433408 310384
rect 433088 310294 433158 310350
rect 433214 310294 433282 310350
rect 433338 310294 433408 310350
rect 433088 310226 433408 310294
rect 433088 310170 433158 310226
rect 433214 310170 433282 310226
rect 433338 310170 433408 310226
rect 433088 310102 433408 310170
rect 433088 310046 433158 310102
rect 433214 310046 433282 310102
rect 433338 310046 433408 310102
rect 433088 309978 433408 310046
rect 433088 309922 433158 309978
rect 433214 309922 433282 309978
rect 433338 309922 433408 309978
rect 433088 309888 433408 309922
rect 435154 310350 435774 327922
rect 435154 310294 435250 310350
rect 435306 310294 435374 310350
rect 435430 310294 435498 310350
rect 435554 310294 435622 310350
rect 435678 310294 435774 310350
rect 435154 310226 435774 310294
rect 435154 310170 435250 310226
rect 435306 310170 435374 310226
rect 435430 310170 435498 310226
rect 435554 310170 435622 310226
rect 435678 310170 435774 310226
rect 435154 310102 435774 310170
rect 435154 310046 435250 310102
rect 435306 310046 435374 310102
rect 435430 310046 435498 310102
rect 435554 310046 435622 310102
rect 435678 310046 435774 310102
rect 435154 309978 435774 310046
rect 435154 309922 435250 309978
rect 435306 309922 435374 309978
rect 435430 309922 435498 309978
rect 435554 309922 435622 309978
rect 435678 309922 435774 309978
rect 420874 298294 420970 298350
rect 421026 298294 421094 298350
rect 421150 298294 421218 298350
rect 421274 298294 421342 298350
rect 421398 298294 421494 298350
rect 420874 298226 421494 298294
rect 420874 298170 420970 298226
rect 421026 298170 421094 298226
rect 421150 298170 421218 298226
rect 421274 298170 421342 298226
rect 421398 298170 421494 298226
rect 420874 298102 421494 298170
rect 420874 298046 420970 298102
rect 421026 298046 421094 298102
rect 421150 298046 421218 298102
rect 421274 298046 421342 298102
rect 421398 298046 421494 298102
rect 420874 297978 421494 298046
rect 420874 297922 420970 297978
rect 421026 297922 421094 297978
rect 421150 297922 421218 297978
rect 421274 297922 421342 297978
rect 421398 297922 421494 297978
rect 402874 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 403494 280350
rect 402874 280226 403494 280294
rect 402874 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 403494 280226
rect 402874 280102 403494 280170
rect 402874 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 403494 280102
rect 402874 279978 403494 280046
rect 402874 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 403494 279978
rect 399154 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 399774 274350
rect 399154 274226 399774 274294
rect 399154 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 399774 274226
rect 399154 274102 399774 274170
rect 399154 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 399774 274102
rect 399154 273978 399774 274046
rect 399154 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 399774 273978
rect 384874 262294 384970 262350
rect 385026 262294 385094 262350
rect 385150 262294 385218 262350
rect 385274 262294 385342 262350
rect 385398 262294 385494 262350
rect 384874 262226 385494 262294
rect 384874 262170 384970 262226
rect 385026 262170 385094 262226
rect 385150 262170 385218 262226
rect 385274 262170 385342 262226
rect 385398 262170 385494 262226
rect 384874 262102 385494 262170
rect 384874 262046 384970 262102
rect 385026 262046 385094 262102
rect 385150 262046 385218 262102
rect 385274 262046 385342 262102
rect 385398 262046 385494 262102
rect 384874 261978 385494 262046
rect 384874 261922 384970 261978
rect 385026 261922 385094 261978
rect 385150 261922 385218 261978
rect 385274 261922 385342 261978
rect 385398 261922 385494 261978
rect 384874 244350 385494 261922
rect 387008 262350 387328 262384
rect 387008 262294 387078 262350
rect 387134 262294 387202 262350
rect 387258 262294 387328 262350
rect 387008 262226 387328 262294
rect 387008 262170 387078 262226
rect 387134 262170 387202 262226
rect 387258 262170 387328 262226
rect 387008 262102 387328 262170
rect 387008 262046 387078 262102
rect 387134 262046 387202 262102
rect 387258 262046 387328 262102
rect 387008 261978 387328 262046
rect 387008 261922 387078 261978
rect 387134 261922 387202 261978
rect 387258 261922 387328 261978
rect 387008 261888 387328 261922
rect 399154 256350 399774 273922
rect 402368 274350 402688 274384
rect 402368 274294 402438 274350
rect 402494 274294 402562 274350
rect 402618 274294 402688 274350
rect 402368 274226 402688 274294
rect 402368 274170 402438 274226
rect 402494 274170 402562 274226
rect 402618 274170 402688 274226
rect 402368 274102 402688 274170
rect 402368 274046 402438 274102
rect 402494 274046 402562 274102
rect 402618 274046 402688 274102
rect 402368 273978 402688 274046
rect 402368 273922 402438 273978
rect 402494 273922 402562 273978
rect 402618 273922 402688 273978
rect 402368 273888 402688 273922
rect 402874 262350 403494 279922
rect 417728 280350 418048 280384
rect 417728 280294 417798 280350
rect 417854 280294 417922 280350
rect 417978 280294 418048 280350
rect 417728 280226 418048 280294
rect 417728 280170 417798 280226
rect 417854 280170 417922 280226
rect 417978 280170 418048 280226
rect 417728 280102 418048 280170
rect 417728 280046 417798 280102
rect 417854 280046 417922 280102
rect 417978 280046 418048 280102
rect 417728 279978 418048 280046
rect 417728 279922 417798 279978
rect 417854 279922 417922 279978
rect 417978 279922 418048 279978
rect 417728 279888 418048 279922
rect 420874 280350 421494 297922
rect 433088 292350 433408 292384
rect 433088 292294 433158 292350
rect 433214 292294 433282 292350
rect 433338 292294 433408 292350
rect 433088 292226 433408 292294
rect 433088 292170 433158 292226
rect 433214 292170 433282 292226
rect 433338 292170 433408 292226
rect 433088 292102 433408 292170
rect 433088 292046 433158 292102
rect 433214 292046 433282 292102
rect 433338 292046 433408 292102
rect 433088 291978 433408 292046
rect 433088 291922 433158 291978
rect 433214 291922 433282 291978
rect 433338 291922 433408 291978
rect 433088 291888 433408 291922
rect 435154 292350 435774 309922
rect 435154 292294 435250 292350
rect 435306 292294 435374 292350
rect 435430 292294 435498 292350
rect 435554 292294 435622 292350
rect 435678 292294 435774 292350
rect 435154 292226 435774 292294
rect 435154 292170 435250 292226
rect 435306 292170 435374 292226
rect 435430 292170 435498 292226
rect 435554 292170 435622 292226
rect 435678 292170 435774 292226
rect 435154 292102 435774 292170
rect 435154 292046 435250 292102
rect 435306 292046 435374 292102
rect 435430 292046 435498 292102
rect 435554 292046 435622 292102
rect 435678 292046 435774 292102
rect 435154 291978 435774 292046
rect 435154 291922 435250 291978
rect 435306 291922 435374 291978
rect 435430 291922 435498 291978
rect 435554 291922 435622 291978
rect 435678 291922 435774 291978
rect 420874 280294 420970 280350
rect 421026 280294 421094 280350
rect 421150 280294 421218 280350
rect 421274 280294 421342 280350
rect 421398 280294 421494 280350
rect 420874 280226 421494 280294
rect 420874 280170 420970 280226
rect 421026 280170 421094 280226
rect 421150 280170 421218 280226
rect 421274 280170 421342 280226
rect 421398 280170 421494 280226
rect 420874 280102 421494 280170
rect 420874 280046 420970 280102
rect 421026 280046 421094 280102
rect 421150 280046 421218 280102
rect 421274 280046 421342 280102
rect 421398 280046 421494 280102
rect 420874 279978 421494 280046
rect 420874 279922 420970 279978
rect 421026 279922 421094 279978
rect 421150 279922 421218 279978
rect 421274 279922 421342 279978
rect 421398 279922 421494 279978
rect 402874 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 403494 262350
rect 402874 262226 403494 262294
rect 402874 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 403494 262226
rect 402874 262102 403494 262170
rect 402874 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 403494 262102
rect 402874 261978 403494 262046
rect 402874 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 403494 261978
rect 399154 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 399774 256350
rect 399154 256226 399774 256294
rect 399154 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 399774 256226
rect 399154 256102 399774 256170
rect 399154 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 399774 256102
rect 399154 255978 399774 256046
rect 399154 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 399774 255978
rect 384874 244294 384970 244350
rect 385026 244294 385094 244350
rect 385150 244294 385218 244350
rect 385274 244294 385342 244350
rect 385398 244294 385494 244350
rect 384874 244226 385494 244294
rect 384874 244170 384970 244226
rect 385026 244170 385094 244226
rect 385150 244170 385218 244226
rect 385274 244170 385342 244226
rect 385398 244170 385494 244226
rect 384874 244102 385494 244170
rect 384874 244046 384970 244102
rect 385026 244046 385094 244102
rect 385150 244046 385218 244102
rect 385274 244046 385342 244102
rect 385398 244046 385494 244102
rect 384874 243978 385494 244046
rect 384874 243922 384970 243978
rect 385026 243922 385094 243978
rect 385150 243922 385218 243978
rect 385274 243922 385342 243978
rect 385398 243922 385494 243978
rect 384874 226350 385494 243922
rect 387008 244350 387328 244384
rect 387008 244294 387078 244350
rect 387134 244294 387202 244350
rect 387258 244294 387328 244350
rect 387008 244226 387328 244294
rect 387008 244170 387078 244226
rect 387134 244170 387202 244226
rect 387258 244170 387328 244226
rect 387008 244102 387328 244170
rect 387008 244046 387078 244102
rect 387134 244046 387202 244102
rect 387258 244046 387328 244102
rect 387008 243978 387328 244046
rect 387008 243922 387078 243978
rect 387134 243922 387202 243978
rect 387258 243922 387328 243978
rect 387008 243888 387328 243922
rect 399154 238350 399774 255922
rect 402368 256350 402688 256384
rect 402368 256294 402438 256350
rect 402494 256294 402562 256350
rect 402618 256294 402688 256350
rect 402368 256226 402688 256294
rect 402368 256170 402438 256226
rect 402494 256170 402562 256226
rect 402618 256170 402688 256226
rect 402368 256102 402688 256170
rect 402368 256046 402438 256102
rect 402494 256046 402562 256102
rect 402618 256046 402688 256102
rect 402368 255978 402688 256046
rect 402368 255922 402438 255978
rect 402494 255922 402562 255978
rect 402618 255922 402688 255978
rect 402368 255888 402688 255922
rect 402874 244350 403494 261922
rect 417728 262350 418048 262384
rect 417728 262294 417798 262350
rect 417854 262294 417922 262350
rect 417978 262294 418048 262350
rect 417728 262226 418048 262294
rect 417728 262170 417798 262226
rect 417854 262170 417922 262226
rect 417978 262170 418048 262226
rect 417728 262102 418048 262170
rect 417728 262046 417798 262102
rect 417854 262046 417922 262102
rect 417978 262046 418048 262102
rect 417728 261978 418048 262046
rect 417728 261922 417798 261978
rect 417854 261922 417922 261978
rect 417978 261922 418048 261978
rect 417728 261888 418048 261922
rect 420874 262350 421494 279922
rect 433088 274350 433408 274384
rect 433088 274294 433158 274350
rect 433214 274294 433282 274350
rect 433338 274294 433408 274350
rect 433088 274226 433408 274294
rect 433088 274170 433158 274226
rect 433214 274170 433282 274226
rect 433338 274170 433408 274226
rect 433088 274102 433408 274170
rect 433088 274046 433158 274102
rect 433214 274046 433282 274102
rect 433338 274046 433408 274102
rect 433088 273978 433408 274046
rect 433088 273922 433158 273978
rect 433214 273922 433282 273978
rect 433338 273922 433408 273978
rect 433088 273888 433408 273922
rect 435154 274350 435774 291922
rect 435154 274294 435250 274350
rect 435306 274294 435374 274350
rect 435430 274294 435498 274350
rect 435554 274294 435622 274350
rect 435678 274294 435774 274350
rect 435154 274226 435774 274294
rect 435154 274170 435250 274226
rect 435306 274170 435374 274226
rect 435430 274170 435498 274226
rect 435554 274170 435622 274226
rect 435678 274170 435774 274226
rect 435154 274102 435774 274170
rect 435154 274046 435250 274102
rect 435306 274046 435374 274102
rect 435430 274046 435498 274102
rect 435554 274046 435622 274102
rect 435678 274046 435774 274102
rect 435154 273978 435774 274046
rect 435154 273922 435250 273978
rect 435306 273922 435374 273978
rect 435430 273922 435498 273978
rect 435554 273922 435622 273978
rect 435678 273922 435774 273978
rect 420874 262294 420970 262350
rect 421026 262294 421094 262350
rect 421150 262294 421218 262350
rect 421274 262294 421342 262350
rect 421398 262294 421494 262350
rect 420874 262226 421494 262294
rect 420874 262170 420970 262226
rect 421026 262170 421094 262226
rect 421150 262170 421218 262226
rect 421274 262170 421342 262226
rect 421398 262170 421494 262226
rect 420874 262102 421494 262170
rect 420874 262046 420970 262102
rect 421026 262046 421094 262102
rect 421150 262046 421218 262102
rect 421274 262046 421342 262102
rect 421398 262046 421494 262102
rect 420874 261978 421494 262046
rect 420874 261922 420970 261978
rect 421026 261922 421094 261978
rect 421150 261922 421218 261978
rect 421274 261922 421342 261978
rect 421398 261922 421494 261978
rect 402874 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 403494 244350
rect 402874 244226 403494 244294
rect 402874 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 403494 244226
rect 402874 244102 403494 244170
rect 402874 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 403494 244102
rect 402874 243978 403494 244046
rect 402874 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 403494 243978
rect 399154 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 399774 238350
rect 399154 238226 399774 238294
rect 399154 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 399774 238226
rect 399154 238102 399774 238170
rect 399154 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 399774 238102
rect 399154 237978 399774 238046
rect 399154 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 399774 237978
rect 384874 226294 384970 226350
rect 385026 226294 385094 226350
rect 385150 226294 385218 226350
rect 385274 226294 385342 226350
rect 385398 226294 385494 226350
rect 384874 226226 385494 226294
rect 384874 226170 384970 226226
rect 385026 226170 385094 226226
rect 385150 226170 385218 226226
rect 385274 226170 385342 226226
rect 385398 226170 385494 226226
rect 384874 226102 385494 226170
rect 384874 226046 384970 226102
rect 385026 226046 385094 226102
rect 385150 226046 385218 226102
rect 385274 226046 385342 226102
rect 385398 226046 385494 226102
rect 384874 225978 385494 226046
rect 384874 225922 384970 225978
rect 385026 225922 385094 225978
rect 385150 225922 385218 225978
rect 385274 225922 385342 225978
rect 385398 225922 385494 225978
rect 384874 208350 385494 225922
rect 387008 226350 387328 226384
rect 387008 226294 387078 226350
rect 387134 226294 387202 226350
rect 387258 226294 387328 226350
rect 387008 226226 387328 226294
rect 387008 226170 387078 226226
rect 387134 226170 387202 226226
rect 387258 226170 387328 226226
rect 387008 226102 387328 226170
rect 387008 226046 387078 226102
rect 387134 226046 387202 226102
rect 387258 226046 387328 226102
rect 387008 225978 387328 226046
rect 387008 225922 387078 225978
rect 387134 225922 387202 225978
rect 387258 225922 387328 225978
rect 387008 225888 387328 225922
rect 399154 220350 399774 237922
rect 402368 238350 402688 238384
rect 402368 238294 402438 238350
rect 402494 238294 402562 238350
rect 402618 238294 402688 238350
rect 402368 238226 402688 238294
rect 402368 238170 402438 238226
rect 402494 238170 402562 238226
rect 402618 238170 402688 238226
rect 402368 238102 402688 238170
rect 402368 238046 402438 238102
rect 402494 238046 402562 238102
rect 402618 238046 402688 238102
rect 402368 237978 402688 238046
rect 402368 237922 402438 237978
rect 402494 237922 402562 237978
rect 402618 237922 402688 237978
rect 402368 237888 402688 237922
rect 402874 226350 403494 243922
rect 417728 244350 418048 244384
rect 417728 244294 417798 244350
rect 417854 244294 417922 244350
rect 417978 244294 418048 244350
rect 417728 244226 418048 244294
rect 417728 244170 417798 244226
rect 417854 244170 417922 244226
rect 417978 244170 418048 244226
rect 417728 244102 418048 244170
rect 417728 244046 417798 244102
rect 417854 244046 417922 244102
rect 417978 244046 418048 244102
rect 417728 243978 418048 244046
rect 417728 243922 417798 243978
rect 417854 243922 417922 243978
rect 417978 243922 418048 243978
rect 417728 243888 418048 243922
rect 420874 244350 421494 261922
rect 433088 256350 433408 256384
rect 433088 256294 433158 256350
rect 433214 256294 433282 256350
rect 433338 256294 433408 256350
rect 433088 256226 433408 256294
rect 433088 256170 433158 256226
rect 433214 256170 433282 256226
rect 433338 256170 433408 256226
rect 433088 256102 433408 256170
rect 433088 256046 433158 256102
rect 433214 256046 433282 256102
rect 433338 256046 433408 256102
rect 433088 255978 433408 256046
rect 433088 255922 433158 255978
rect 433214 255922 433282 255978
rect 433338 255922 433408 255978
rect 433088 255888 433408 255922
rect 435154 256350 435774 273922
rect 435154 256294 435250 256350
rect 435306 256294 435374 256350
rect 435430 256294 435498 256350
rect 435554 256294 435622 256350
rect 435678 256294 435774 256350
rect 435154 256226 435774 256294
rect 435154 256170 435250 256226
rect 435306 256170 435374 256226
rect 435430 256170 435498 256226
rect 435554 256170 435622 256226
rect 435678 256170 435774 256226
rect 435154 256102 435774 256170
rect 435154 256046 435250 256102
rect 435306 256046 435374 256102
rect 435430 256046 435498 256102
rect 435554 256046 435622 256102
rect 435678 256046 435774 256102
rect 435154 255978 435774 256046
rect 435154 255922 435250 255978
rect 435306 255922 435374 255978
rect 435430 255922 435498 255978
rect 435554 255922 435622 255978
rect 435678 255922 435774 255978
rect 420874 244294 420970 244350
rect 421026 244294 421094 244350
rect 421150 244294 421218 244350
rect 421274 244294 421342 244350
rect 421398 244294 421494 244350
rect 420874 244226 421494 244294
rect 420874 244170 420970 244226
rect 421026 244170 421094 244226
rect 421150 244170 421218 244226
rect 421274 244170 421342 244226
rect 421398 244170 421494 244226
rect 420874 244102 421494 244170
rect 420874 244046 420970 244102
rect 421026 244046 421094 244102
rect 421150 244046 421218 244102
rect 421274 244046 421342 244102
rect 421398 244046 421494 244102
rect 420874 243978 421494 244046
rect 420874 243922 420970 243978
rect 421026 243922 421094 243978
rect 421150 243922 421218 243978
rect 421274 243922 421342 243978
rect 421398 243922 421494 243978
rect 402874 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 403494 226350
rect 402874 226226 403494 226294
rect 402874 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 403494 226226
rect 402874 226102 403494 226170
rect 402874 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 403494 226102
rect 402874 225978 403494 226046
rect 402874 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 403494 225978
rect 399154 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 399774 220350
rect 399154 220226 399774 220294
rect 399154 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 399774 220226
rect 399154 220102 399774 220170
rect 399154 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 399774 220102
rect 399154 219978 399774 220046
rect 399154 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 399774 219978
rect 384874 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 385494 208350
rect 384874 208226 385494 208294
rect 384874 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 385494 208226
rect 384874 208102 385494 208170
rect 384874 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 385494 208102
rect 384874 207978 385494 208046
rect 384874 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 385494 207978
rect 384874 190350 385494 207922
rect 387008 208350 387328 208384
rect 387008 208294 387078 208350
rect 387134 208294 387202 208350
rect 387258 208294 387328 208350
rect 387008 208226 387328 208294
rect 387008 208170 387078 208226
rect 387134 208170 387202 208226
rect 387258 208170 387328 208226
rect 387008 208102 387328 208170
rect 387008 208046 387078 208102
rect 387134 208046 387202 208102
rect 387258 208046 387328 208102
rect 387008 207978 387328 208046
rect 387008 207922 387078 207978
rect 387134 207922 387202 207978
rect 387258 207922 387328 207978
rect 387008 207888 387328 207922
rect 399154 202350 399774 219922
rect 402368 220350 402688 220384
rect 402368 220294 402438 220350
rect 402494 220294 402562 220350
rect 402618 220294 402688 220350
rect 402368 220226 402688 220294
rect 402368 220170 402438 220226
rect 402494 220170 402562 220226
rect 402618 220170 402688 220226
rect 402368 220102 402688 220170
rect 402368 220046 402438 220102
rect 402494 220046 402562 220102
rect 402618 220046 402688 220102
rect 402368 219978 402688 220046
rect 402368 219922 402438 219978
rect 402494 219922 402562 219978
rect 402618 219922 402688 219978
rect 402368 219888 402688 219922
rect 402874 208350 403494 225922
rect 417728 226350 418048 226384
rect 417728 226294 417798 226350
rect 417854 226294 417922 226350
rect 417978 226294 418048 226350
rect 417728 226226 418048 226294
rect 417728 226170 417798 226226
rect 417854 226170 417922 226226
rect 417978 226170 418048 226226
rect 417728 226102 418048 226170
rect 417728 226046 417798 226102
rect 417854 226046 417922 226102
rect 417978 226046 418048 226102
rect 417728 225978 418048 226046
rect 417728 225922 417798 225978
rect 417854 225922 417922 225978
rect 417978 225922 418048 225978
rect 417728 225888 418048 225922
rect 420874 226350 421494 243922
rect 433088 238350 433408 238384
rect 433088 238294 433158 238350
rect 433214 238294 433282 238350
rect 433338 238294 433408 238350
rect 433088 238226 433408 238294
rect 433088 238170 433158 238226
rect 433214 238170 433282 238226
rect 433338 238170 433408 238226
rect 433088 238102 433408 238170
rect 433088 238046 433158 238102
rect 433214 238046 433282 238102
rect 433338 238046 433408 238102
rect 433088 237978 433408 238046
rect 433088 237922 433158 237978
rect 433214 237922 433282 237978
rect 433338 237922 433408 237978
rect 433088 237888 433408 237922
rect 435154 238350 435774 255922
rect 435154 238294 435250 238350
rect 435306 238294 435374 238350
rect 435430 238294 435498 238350
rect 435554 238294 435622 238350
rect 435678 238294 435774 238350
rect 435154 238226 435774 238294
rect 435154 238170 435250 238226
rect 435306 238170 435374 238226
rect 435430 238170 435498 238226
rect 435554 238170 435622 238226
rect 435678 238170 435774 238226
rect 435154 238102 435774 238170
rect 435154 238046 435250 238102
rect 435306 238046 435374 238102
rect 435430 238046 435498 238102
rect 435554 238046 435622 238102
rect 435678 238046 435774 238102
rect 435154 237978 435774 238046
rect 435154 237922 435250 237978
rect 435306 237922 435374 237978
rect 435430 237922 435498 237978
rect 435554 237922 435622 237978
rect 435678 237922 435774 237978
rect 420874 226294 420970 226350
rect 421026 226294 421094 226350
rect 421150 226294 421218 226350
rect 421274 226294 421342 226350
rect 421398 226294 421494 226350
rect 420874 226226 421494 226294
rect 420874 226170 420970 226226
rect 421026 226170 421094 226226
rect 421150 226170 421218 226226
rect 421274 226170 421342 226226
rect 421398 226170 421494 226226
rect 420874 226102 421494 226170
rect 420874 226046 420970 226102
rect 421026 226046 421094 226102
rect 421150 226046 421218 226102
rect 421274 226046 421342 226102
rect 421398 226046 421494 226102
rect 420874 225978 421494 226046
rect 420874 225922 420970 225978
rect 421026 225922 421094 225978
rect 421150 225922 421218 225978
rect 421274 225922 421342 225978
rect 421398 225922 421494 225978
rect 402874 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 403494 208350
rect 402874 208226 403494 208294
rect 402874 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 403494 208226
rect 402874 208102 403494 208170
rect 402874 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 403494 208102
rect 402874 207978 403494 208046
rect 402874 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 403494 207978
rect 399154 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 399774 202350
rect 399154 202226 399774 202294
rect 399154 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 399774 202226
rect 399154 202102 399774 202170
rect 399154 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 399774 202102
rect 399154 201978 399774 202046
rect 399154 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 399774 201978
rect 384874 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 385494 190350
rect 384874 190226 385494 190294
rect 384874 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 385494 190226
rect 384874 190102 385494 190170
rect 384874 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 385494 190102
rect 384874 189978 385494 190046
rect 384874 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 385494 189978
rect 384874 172350 385494 189922
rect 387008 190350 387328 190384
rect 387008 190294 387078 190350
rect 387134 190294 387202 190350
rect 387258 190294 387328 190350
rect 387008 190226 387328 190294
rect 387008 190170 387078 190226
rect 387134 190170 387202 190226
rect 387258 190170 387328 190226
rect 387008 190102 387328 190170
rect 387008 190046 387078 190102
rect 387134 190046 387202 190102
rect 387258 190046 387328 190102
rect 387008 189978 387328 190046
rect 387008 189922 387078 189978
rect 387134 189922 387202 189978
rect 387258 189922 387328 189978
rect 387008 189888 387328 189922
rect 399154 184350 399774 201922
rect 402368 202350 402688 202384
rect 402368 202294 402438 202350
rect 402494 202294 402562 202350
rect 402618 202294 402688 202350
rect 402368 202226 402688 202294
rect 402368 202170 402438 202226
rect 402494 202170 402562 202226
rect 402618 202170 402688 202226
rect 402368 202102 402688 202170
rect 402368 202046 402438 202102
rect 402494 202046 402562 202102
rect 402618 202046 402688 202102
rect 402368 201978 402688 202046
rect 402368 201922 402438 201978
rect 402494 201922 402562 201978
rect 402618 201922 402688 201978
rect 402368 201888 402688 201922
rect 402874 190350 403494 207922
rect 417728 208350 418048 208384
rect 417728 208294 417798 208350
rect 417854 208294 417922 208350
rect 417978 208294 418048 208350
rect 417728 208226 418048 208294
rect 417728 208170 417798 208226
rect 417854 208170 417922 208226
rect 417978 208170 418048 208226
rect 417728 208102 418048 208170
rect 417728 208046 417798 208102
rect 417854 208046 417922 208102
rect 417978 208046 418048 208102
rect 417728 207978 418048 208046
rect 417728 207922 417798 207978
rect 417854 207922 417922 207978
rect 417978 207922 418048 207978
rect 417728 207888 418048 207922
rect 420874 208350 421494 225922
rect 433088 220350 433408 220384
rect 433088 220294 433158 220350
rect 433214 220294 433282 220350
rect 433338 220294 433408 220350
rect 433088 220226 433408 220294
rect 433088 220170 433158 220226
rect 433214 220170 433282 220226
rect 433338 220170 433408 220226
rect 433088 220102 433408 220170
rect 433088 220046 433158 220102
rect 433214 220046 433282 220102
rect 433338 220046 433408 220102
rect 433088 219978 433408 220046
rect 433088 219922 433158 219978
rect 433214 219922 433282 219978
rect 433338 219922 433408 219978
rect 433088 219888 433408 219922
rect 435154 220350 435774 237922
rect 435154 220294 435250 220350
rect 435306 220294 435374 220350
rect 435430 220294 435498 220350
rect 435554 220294 435622 220350
rect 435678 220294 435774 220350
rect 435154 220226 435774 220294
rect 435154 220170 435250 220226
rect 435306 220170 435374 220226
rect 435430 220170 435498 220226
rect 435554 220170 435622 220226
rect 435678 220170 435774 220226
rect 435154 220102 435774 220170
rect 435154 220046 435250 220102
rect 435306 220046 435374 220102
rect 435430 220046 435498 220102
rect 435554 220046 435622 220102
rect 435678 220046 435774 220102
rect 435154 219978 435774 220046
rect 435154 219922 435250 219978
rect 435306 219922 435374 219978
rect 435430 219922 435498 219978
rect 435554 219922 435622 219978
rect 435678 219922 435774 219978
rect 420874 208294 420970 208350
rect 421026 208294 421094 208350
rect 421150 208294 421218 208350
rect 421274 208294 421342 208350
rect 421398 208294 421494 208350
rect 420874 208226 421494 208294
rect 420874 208170 420970 208226
rect 421026 208170 421094 208226
rect 421150 208170 421218 208226
rect 421274 208170 421342 208226
rect 421398 208170 421494 208226
rect 420874 208102 421494 208170
rect 420874 208046 420970 208102
rect 421026 208046 421094 208102
rect 421150 208046 421218 208102
rect 421274 208046 421342 208102
rect 421398 208046 421494 208102
rect 420874 207978 421494 208046
rect 420874 207922 420970 207978
rect 421026 207922 421094 207978
rect 421150 207922 421218 207978
rect 421274 207922 421342 207978
rect 421398 207922 421494 207978
rect 402874 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 403494 190350
rect 402874 190226 403494 190294
rect 402874 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 403494 190226
rect 402874 190102 403494 190170
rect 402874 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 403494 190102
rect 402874 189978 403494 190046
rect 402874 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 403494 189978
rect 399154 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 399774 184350
rect 399154 184226 399774 184294
rect 399154 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 399774 184226
rect 399154 184102 399774 184170
rect 399154 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 399774 184102
rect 399154 183978 399774 184046
rect 399154 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 399774 183978
rect 384874 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 385494 172350
rect 384874 172226 385494 172294
rect 384874 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 385494 172226
rect 384874 172102 385494 172170
rect 384874 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 385494 172102
rect 384874 171978 385494 172046
rect 384874 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 385494 171978
rect 384874 154350 385494 171922
rect 387008 172350 387328 172384
rect 387008 172294 387078 172350
rect 387134 172294 387202 172350
rect 387258 172294 387328 172350
rect 387008 172226 387328 172294
rect 387008 172170 387078 172226
rect 387134 172170 387202 172226
rect 387258 172170 387328 172226
rect 387008 172102 387328 172170
rect 387008 172046 387078 172102
rect 387134 172046 387202 172102
rect 387258 172046 387328 172102
rect 387008 171978 387328 172046
rect 387008 171922 387078 171978
rect 387134 171922 387202 171978
rect 387258 171922 387328 171978
rect 387008 171888 387328 171922
rect 399154 166350 399774 183922
rect 402368 184350 402688 184384
rect 402368 184294 402438 184350
rect 402494 184294 402562 184350
rect 402618 184294 402688 184350
rect 402368 184226 402688 184294
rect 402368 184170 402438 184226
rect 402494 184170 402562 184226
rect 402618 184170 402688 184226
rect 402368 184102 402688 184170
rect 402368 184046 402438 184102
rect 402494 184046 402562 184102
rect 402618 184046 402688 184102
rect 402368 183978 402688 184046
rect 402368 183922 402438 183978
rect 402494 183922 402562 183978
rect 402618 183922 402688 183978
rect 402368 183888 402688 183922
rect 402874 172350 403494 189922
rect 417728 190350 418048 190384
rect 417728 190294 417798 190350
rect 417854 190294 417922 190350
rect 417978 190294 418048 190350
rect 417728 190226 418048 190294
rect 417728 190170 417798 190226
rect 417854 190170 417922 190226
rect 417978 190170 418048 190226
rect 417728 190102 418048 190170
rect 417728 190046 417798 190102
rect 417854 190046 417922 190102
rect 417978 190046 418048 190102
rect 417728 189978 418048 190046
rect 417728 189922 417798 189978
rect 417854 189922 417922 189978
rect 417978 189922 418048 189978
rect 417728 189888 418048 189922
rect 420874 190350 421494 207922
rect 433088 202350 433408 202384
rect 433088 202294 433158 202350
rect 433214 202294 433282 202350
rect 433338 202294 433408 202350
rect 433088 202226 433408 202294
rect 433088 202170 433158 202226
rect 433214 202170 433282 202226
rect 433338 202170 433408 202226
rect 433088 202102 433408 202170
rect 433088 202046 433158 202102
rect 433214 202046 433282 202102
rect 433338 202046 433408 202102
rect 433088 201978 433408 202046
rect 433088 201922 433158 201978
rect 433214 201922 433282 201978
rect 433338 201922 433408 201978
rect 433088 201888 433408 201922
rect 435154 202350 435774 219922
rect 435154 202294 435250 202350
rect 435306 202294 435374 202350
rect 435430 202294 435498 202350
rect 435554 202294 435622 202350
rect 435678 202294 435774 202350
rect 435154 202226 435774 202294
rect 435154 202170 435250 202226
rect 435306 202170 435374 202226
rect 435430 202170 435498 202226
rect 435554 202170 435622 202226
rect 435678 202170 435774 202226
rect 435154 202102 435774 202170
rect 435154 202046 435250 202102
rect 435306 202046 435374 202102
rect 435430 202046 435498 202102
rect 435554 202046 435622 202102
rect 435678 202046 435774 202102
rect 435154 201978 435774 202046
rect 435154 201922 435250 201978
rect 435306 201922 435374 201978
rect 435430 201922 435498 201978
rect 435554 201922 435622 201978
rect 435678 201922 435774 201978
rect 420874 190294 420970 190350
rect 421026 190294 421094 190350
rect 421150 190294 421218 190350
rect 421274 190294 421342 190350
rect 421398 190294 421494 190350
rect 420874 190226 421494 190294
rect 420874 190170 420970 190226
rect 421026 190170 421094 190226
rect 421150 190170 421218 190226
rect 421274 190170 421342 190226
rect 421398 190170 421494 190226
rect 420874 190102 421494 190170
rect 420874 190046 420970 190102
rect 421026 190046 421094 190102
rect 421150 190046 421218 190102
rect 421274 190046 421342 190102
rect 421398 190046 421494 190102
rect 420874 189978 421494 190046
rect 420874 189922 420970 189978
rect 421026 189922 421094 189978
rect 421150 189922 421218 189978
rect 421274 189922 421342 189978
rect 421398 189922 421494 189978
rect 402874 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 403494 172350
rect 402874 172226 403494 172294
rect 402874 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 403494 172226
rect 402874 172102 403494 172170
rect 402874 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 403494 172102
rect 402874 171978 403494 172046
rect 402874 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 403494 171978
rect 399154 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 399774 166350
rect 399154 166226 399774 166294
rect 399154 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 399774 166226
rect 399154 166102 399774 166170
rect 399154 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 399774 166102
rect 399154 165978 399774 166046
rect 399154 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 399774 165978
rect 384874 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 385494 154350
rect 384874 154226 385494 154294
rect 384874 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 385494 154226
rect 384874 154102 385494 154170
rect 384874 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 385494 154102
rect 384874 153978 385494 154046
rect 384874 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 385494 153978
rect 384874 136350 385494 153922
rect 387008 154350 387328 154384
rect 387008 154294 387078 154350
rect 387134 154294 387202 154350
rect 387258 154294 387328 154350
rect 387008 154226 387328 154294
rect 387008 154170 387078 154226
rect 387134 154170 387202 154226
rect 387258 154170 387328 154226
rect 387008 154102 387328 154170
rect 387008 154046 387078 154102
rect 387134 154046 387202 154102
rect 387258 154046 387328 154102
rect 387008 153978 387328 154046
rect 387008 153922 387078 153978
rect 387134 153922 387202 153978
rect 387258 153922 387328 153978
rect 387008 153888 387328 153922
rect 399154 148350 399774 165922
rect 402368 166350 402688 166384
rect 402368 166294 402438 166350
rect 402494 166294 402562 166350
rect 402618 166294 402688 166350
rect 402368 166226 402688 166294
rect 402368 166170 402438 166226
rect 402494 166170 402562 166226
rect 402618 166170 402688 166226
rect 402368 166102 402688 166170
rect 402368 166046 402438 166102
rect 402494 166046 402562 166102
rect 402618 166046 402688 166102
rect 402368 165978 402688 166046
rect 402368 165922 402438 165978
rect 402494 165922 402562 165978
rect 402618 165922 402688 165978
rect 402368 165888 402688 165922
rect 402874 154350 403494 171922
rect 417728 172350 418048 172384
rect 417728 172294 417798 172350
rect 417854 172294 417922 172350
rect 417978 172294 418048 172350
rect 417728 172226 418048 172294
rect 417728 172170 417798 172226
rect 417854 172170 417922 172226
rect 417978 172170 418048 172226
rect 417728 172102 418048 172170
rect 417728 172046 417798 172102
rect 417854 172046 417922 172102
rect 417978 172046 418048 172102
rect 417728 171978 418048 172046
rect 417728 171922 417798 171978
rect 417854 171922 417922 171978
rect 417978 171922 418048 171978
rect 417728 171888 418048 171922
rect 420874 172350 421494 189922
rect 433088 184350 433408 184384
rect 433088 184294 433158 184350
rect 433214 184294 433282 184350
rect 433338 184294 433408 184350
rect 433088 184226 433408 184294
rect 433088 184170 433158 184226
rect 433214 184170 433282 184226
rect 433338 184170 433408 184226
rect 433088 184102 433408 184170
rect 433088 184046 433158 184102
rect 433214 184046 433282 184102
rect 433338 184046 433408 184102
rect 433088 183978 433408 184046
rect 433088 183922 433158 183978
rect 433214 183922 433282 183978
rect 433338 183922 433408 183978
rect 433088 183888 433408 183922
rect 435154 184350 435774 201922
rect 435154 184294 435250 184350
rect 435306 184294 435374 184350
rect 435430 184294 435498 184350
rect 435554 184294 435622 184350
rect 435678 184294 435774 184350
rect 435154 184226 435774 184294
rect 435154 184170 435250 184226
rect 435306 184170 435374 184226
rect 435430 184170 435498 184226
rect 435554 184170 435622 184226
rect 435678 184170 435774 184226
rect 435154 184102 435774 184170
rect 435154 184046 435250 184102
rect 435306 184046 435374 184102
rect 435430 184046 435498 184102
rect 435554 184046 435622 184102
rect 435678 184046 435774 184102
rect 435154 183978 435774 184046
rect 435154 183922 435250 183978
rect 435306 183922 435374 183978
rect 435430 183922 435498 183978
rect 435554 183922 435622 183978
rect 435678 183922 435774 183978
rect 420874 172294 420970 172350
rect 421026 172294 421094 172350
rect 421150 172294 421218 172350
rect 421274 172294 421342 172350
rect 421398 172294 421494 172350
rect 420874 172226 421494 172294
rect 420874 172170 420970 172226
rect 421026 172170 421094 172226
rect 421150 172170 421218 172226
rect 421274 172170 421342 172226
rect 421398 172170 421494 172226
rect 420874 172102 421494 172170
rect 420874 172046 420970 172102
rect 421026 172046 421094 172102
rect 421150 172046 421218 172102
rect 421274 172046 421342 172102
rect 421398 172046 421494 172102
rect 420874 171978 421494 172046
rect 420874 171922 420970 171978
rect 421026 171922 421094 171978
rect 421150 171922 421218 171978
rect 421274 171922 421342 171978
rect 421398 171922 421494 171978
rect 402874 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 403494 154350
rect 402874 154226 403494 154294
rect 402874 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 403494 154226
rect 402874 154102 403494 154170
rect 402874 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 403494 154102
rect 402874 153978 403494 154046
rect 402874 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 403494 153978
rect 399154 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 399774 148350
rect 399154 148226 399774 148294
rect 399154 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 399774 148226
rect 399154 148102 399774 148170
rect 399154 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 399774 148102
rect 399154 147978 399774 148046
rect 399154 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 399774 147978
rect 384874 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 385494 136350
rect 384874 136226 385494 136294
rect 384874 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 385494 136226
rect 384874 136102 385494 136170
rect 384874 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 385494 136102
rect 384874 135978 385494 136046
rect 384874 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 385494 135978
rect 384874 118350 385494 135922
rect 387008 136350 387328 136384
rect 387008 136294 387078 136350
rect 387134 136294 387202 136350
rect 387258 136294 387328 136350
rect 387008 136226 387328 136294
rect 387008 136170 387078 136226
rect 387134 136170 387202 136226
rect 387258 136170 387328 136226
rect 387008 136102 387328 136170
rect 387008 136046 387078 136102
rect 387134 136046 387202 136102
rect 387258 136046 387328 136102
rect 387008 135978 387328 136046
rect 387008 135922 387078 135978
rect 387134 135922 387202 135978
rect 387258 135922 387328 135978
rect 387008 135888 387328 135922
rect 399154 130350 399774 147922
rect 402368 148350 402688 148384
rect 402368 148294 402438 148350
rect 402494 148294 402562 148350
rect 402618 148294 402688 148350
rect 402368 148226 402688 148294
rect 402368 148170 402438 148226
rect 402494 148170 402562 148226
rect 402618 148170 402688 148226
rect 402368 148102 402688 148170
rect 402368 148046 402438 148102
rect 402494 148046 402562 148102
rect 402618 148046 402688 148102
rect 402368 147978 402688 148046
rect 402368 147922 402438 147978
rect 402494 147922 402562 147978
rect 402618 147922 402688 147978
rect 402368 147888 402688 147922
rect 402874 136350 403494 153922
rect 417728 154350 418048 154384
rect 417728 154294 417798 154350
rect 417854 154294 417922 154350
rect 417978 154294 418048 154350
rect 417728 154226 418048 154294
rect 417728 154170 417798 154226
rect 417854 154170 417922 154226
rect 417978 154170 418048 154226
rect 417728 154102 418048 154170
rect 417728 154046 417798 154102
rect 417854 154046 417922 154102
rect 417978 154046 418048 154102
rect 417728 153978 418048 154046
rect 417728 153922 417798 153978
rect 417854 153922 417922 153978
rect 417978 153922 418048 153978
rect 417728 153888 418048 153922
rect 420874 154350 421494 171922
rect 433088 166350 433408 166384
rect 433088 166294 433158 166350
rect 433214 166294 433282 166350
rect 433338 166294 433408 166350
rect 433088 166226 433408 166294
rect 433088 166170 433158 166226
rect 433214 166170 433282 166226
rect 433338 166170 433408 166226
rect 433088 166102 433408 166170
rect 433088 166046 433158 166102
rect 433214 166046 433282 166102
rect 433338 166046 433408 166102
rect 433088 165978 433408 166046
rect 433088 165922 433158 165978
rect 433214 165922 433282 165978
rect 433338 165922 433408 165978
rect 433088 165888 433408 165922
rect 435154 166350 435774 183922
rect 435154 166294 435250 166350
rect 435306 166294 435374 166350
rect 435430 166294 435498 166350
rect 435554 166294 435622 166350
rect 435678 166294 435774 166350
rect 435154 166226 435774 166294
rect 435154 166170 435250 166226
rect 435306 166170 435374 166226
rect 435430 166170 435498 166226
rect 435554 166170 435622 166226
rect 435678 166170 435774 166226
rect 435154 166102 435774 166170
rect 435154 166046 435250 166102
rect 435306 166046 435374 166102
rect 435430 166046 435498 166102
rect 435554 166046 435622 166102
rect 435678 166046 435774 166102
rect 435154 165978 435774 166046
rect 435154 165922 435250 165978
rect 435306 165922 435374 165978
rect 435430 165922 435498 165978
rect 435554 165922 435622 165978
rect 435678 165922 435774 165978
rect 420874 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 421494 154350
rect 420874 154226 421494 154294
rect 420874 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 421494 154226
rect 420874 154102 421494 154170
rect 420874 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 421494 154102
rect 420874 153978 421494 154046
rect 420874 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 421494 153978
rect 402874 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 403494 136350
rect 402874 136226 403494 136294
rect 402874 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 403494 136226
rect 402874 136102 403494 136170
rect 402874 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 403494 136102
rect 402874 135978 403494 136046
rect 402874 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 403494 135978
rect 399154 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 399774 130350
rect 399154 130226 399774 130294
rect 399154 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 399774 130226
rect 399154 130102 399774 130170
rect 399154 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 399774 130102
rect 399154 129978 399774 130046
rect 399154 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 399774 129978
rect 384874 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 385494 118350
rect 384874 118226 385494 118294
rect 384874 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 385494 118226
rect 384874 118102 385494 118170
rect 384874 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 385494 118102
rect 384874 117978 385494 118046
rect 384874 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 385494 117978
rect 384874 100350 385494 117922
rect 387008 118350 387328 118384
rect 387008 118294 387078 118350
rect 387134 118294 387202 118350
rect 387258 118294 387328 118350
rect 387008 118226 387328 118294
rect 387008 118170 387078 118226
rect 387134 118170 387202 118226
rect 387258 118170 387328 118226
rect 387008 118102 387328 118170
rect 387008 118046 387078 118102
rect 387134 118046 387202 118102
rect 387258 118046 387328 118102
rect 387008 117978 387328 118046
rect 387008 117922 387078 117978
rect 387134 117922 387202 117978
rect 387258 117922 387328 117978
rect 387008 117888 387328 117922
rect 399154 112350 399774 129922
rect 402368 130350 402688 130384
rect 402368 130294 402438 130350
rect 402494 130294 402562 130350
rect 402618 130294 402688 130350
rect 402368 130226 402688 130294
rect 402368 130170 402438 130226
rect 402494 130170 402562 130226
rect 402618 130170 402688 130226
rect 402368 130102 402688 130170
rect 402368 130046 402438 130102
rect 402494 130046 402562 130102
rect 402618 130046 402688 130102
rect 402368 129978 402688 130046
rect 402368 129922 402438 129978
rect 402494 129922 402562 129978
rect 402618 129922 402688 129978
rect 402368 129888 402688 129922
rect 402874 118350 403494 135922
rect 417728 136350 418048 136384
rect 417728 136294 417798 136350
rect 417854 136294 417922 136350
rect 417978 136294 418048 136350
rect 417728 136226 418048 136294
rect 417728 136170 417798 136226
rect 417854 136170 417922 136226
rect 417978 136170 418048 136226
rect 417728 136102 418048 136170
rect 417728 136046 417798 136102
rect 417854 136046 417922 136102
rect 417978 136046 418048 136102
rect 417728 135978 418048 136046
rect 417728 135922 417798 135978
rect 417854 135922 417922 135978
rect 417978 135922 418048 135978
rect 417728 135888 418048 135922
rect 420874 136350 421494 153922
rect 433088 148350 433408 148384
rect 433088 148294 433158 148350
rect 433214 148294 433282 148350
rect 433338 148294 433408 148350
rect 433088 148226 433408 148294
rect 433088 148170 433158 148226
rect 433214 148170 433282 148226
rect 433338 148170 433408 148226
rect 433088 148102 433408 148170
rect 433088 148046 433158 148102
rect 433214 148046 433282 148102
rect 433338 148046 433408 148102
rect 433088 147978 433408 148046
rect 433088 147922 433158 147978
rect 433214 147922 433282 147978
rect 433338 147922 433408 147978
rect 433088 147888 433408 147922
rect 435154 148350 435774 165922
rect 435154 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 435774 148350
rect 435154 148226 435774 148294
rect 435154 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 435774 148226
rect 435154 148102 435774 148170
rect 435154 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 435774 148102
rect 435154 147978 435774 148046
rect 435154 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 435774 147978
rect 420874 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 421494 136350
rect 420874 136226 421494 136294
rect 420874 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 421494 136226
rect 420874 136102 421494 136170
rect 420874 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 421494 136102
rect 420874 135978 421494 136046
rect 420874 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 421494 135978
rect 402874 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 403494 118350
rect 402874 118226 403494 118294
rect 402874 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 403494 118226
rect 402874 118102 403494 118170
rect 402874 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 403494 118102
rect 402874 117978 403494 118046
rect 402874 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 403494 117978
rect 399154 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 399774 112350
rect 399154 112226 399774 112294
rect 399154 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 399774 112226
rect 399154 112102 399774 112170
rect 399154 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 399774 112102
rect 399154 111978 399774 112046
rect 399154 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 399774 111978
rect 384874 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 385494 100350
rect 384874 100226 385494 100294
rect 384874 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 385494 100226
rect 384874 100102 385494 100170
rect 384874 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 385494 100102
rect 384874 99978 385494 100046
rect 384874 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 385494 99978
rect 384874 82350 385494 99922
rect 387008 100350 387328 100384
rect 387008 100294 387078 100350
rect 387134 100294 387202 100350
rect 387258 100294 387328 100350
rect 387008 100226 387328 100294
rect 387008 100170 387078 100226
rect 387134 100170 387202 100226
rect 387258 100170 387328 100226
rect 387008 100102 387328 100170
rect 387008 100046 387078 100102
rect 387134 100046 387202 100102
rect 387258 100046 387328 100102
rect 387008 99978 387328 100046
rect 387008 99922 387078 99978
rect 387134 99922 387202 99978
rect 387258 99922 387328 99978
rect 387008 99888 387328 99922
rect 399154 94350 399774 111922
rect 402368 112350 402688 112384
rect 402368 112294 402438 112350
rect 402494 112294 402562 112350
rect 402618 112294 402688 112350
rect 402368 112226 402688 112294
rect 402368 112170 402438 112226
rect 402494 112170 402562 112226
rect 402618 112170 402688 112226
rect 402368 112102 402688 112170
rect 402368 112046 402438 112102
rect 402494 112046 402562 112102
rect 402618 112046 402688 112102
rect 402368 111978 402688 112046
rect 402368 111922 402438 111978
rect 402494 111922 402562 111978
rect 402618 111922 402688 111978
rect 402368 111888 402688 111922
rect 402874 100350 403494 117922
rect 417728 118350 418048 118384
rect 417728 118294 417798 118350
rect 417854 118294 417922 118350
rect 417978 118294 418048 118350
rect 417728 118226 418048 118294
rect 417728 118170 417798 118226
rect 417854 118170 417922 118226
rect 417978 118170 418048 118226
rect 417728 118102 418048 118170
rect 417728 118046 417798 118102
rect 417854 118046 417922 118102
rect 417978 118046 418048 118102
rect 417728 117978 418048 118046
rect 417728 117922 417798 117978
rect 417854 117922 417922 117978
rect 417978 117922 418048 117978
rect 417728 117888 418048 117922
rect 420874 118350 421494 135922
rect 433088 130350 433408 130384
rect 433088 130294 433158 130350
rect 433214 130294 433282 130350
rect 433338 130294 433408 130350
rect 433088 130226 433408 130294
rect 433088 130170 433158 130226
rect 433214 130170 433282 130226
rect 433338 130170 433408 130226
rect 433088 130102 433408 130170
rect 433088 130046 433158 130102
rect 433214 130046 433282 130102
rect 433338 130046 433408 130102
rect 433088 129978 433408 130046
rect 433088 129922 433158 129978
rect 433214 129922 433282 129978
rect 433338 129922 433408 129978
rect 433088 129888 433408 129922
rect 435154 130350 435774 147922
rect 435154 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 435774 130350
rect 435154 130226 435774 130294
rect 435154 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 435774 130226
rect 435154 130102 435774 130170
rect 435154 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 435774 130102
rect 435154 129978 435774 130046
rect 435154 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 435774 129978
rect 420874 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 421494 118350
rect 420874 118226 421494 118294
rect 420874 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 421494 118226
rect 420874 118102 421494 118170
rect 420874 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 421494 118102
rect 420874 117978 421494 118046
rect 420874 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 421494 117978
rect 402874 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 403494 100350
rect 402874 100226 403494 100294
rect 402874 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 403494 100226
rect 402874 100102 403494 100170
rect 402874 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 403494 100102
rect 402874 99978 403494 100046
rect 402874 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 403494 99978
rect 399154 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 399774 94350
rect 399154 94226 399774 94294
rect 399154 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 399774 94226
rect 399154 94102 399774 94170
rect 399154 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 399774 94102
rect 399154 93978 399774 94046
rect 399154 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 399774 93978
rect 384874 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 385494 82350
rect 384874 82226 385494 82294
rect 384874 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 385494 82226
rect 384874 82102 385494 82170
rect 384874 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 385494 82102
rect 384874 81978 385494 82046
rect 384874 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 385494 81978
rect 384874 64350 385494 81922
rect 387008 82350 387328 82384
rect 387008 82294 387078 82350
rect 387134 82294 387202 82350
rect 387258 82294 387328 82350
rect 387008 82226 387328 82294
rect 387008 82170 387078 82226
rect 387134 82170 387202 82226
rect 387258 82170 387328 82226
rect 387008 82102 387328 82170
rect 387008 82046 387078 82102
rect 387134 82046 387202 82102
rect 387258 82046 387328 82102
rect 387008 81978 387328 82046
rect 387008 81922 387078 81978
rect 387134 81922 387202 81978
rect 387258 81922 387328 81978
rect 387008 81888 387328 81922
rect 399154 76350 399774 93922
rect 402368 94350 402688 94384
rect 402368 94294 402438 94350
rect 402494 94294 402562 94350
rect 402618 94294 402688 94350
rect 402368 94226 402688 94294
rect 402368 94170 402438 94226
rect 402494 94170 402562 94226
rect 402618 94170 402688 94226
rect 402368 94102 402688 94170
rect 402368 94046 402438 94102
rect 402494 94046 402562 94102
rect 402618 94046 402688 94102
rect 402368 93978 402688 94046
rect 402368 93922 402438 93978
rect 402494 93922 402562 93978
rect 402618 93922 402688 93978
rect 402368 93888 402688 93922
rect 402874 82350 403494 99922
rect 417728 100350 418048 100384
rect 417728 100294 417798 100350
rect 417854 100294 417922 100350
rect 417978 100294 418048 100350
rect 417728 100226 418048 100294
rect 417728 100170 417798 100226
rect 417854 100170 417922 100226
rect 417978 100170 418048 100226
rect 417728 100102 418048 100170
rect 417728 100046 417798 100102
rect 417854 100046 417922 100102
rect 417978 100046 418048 100102
rect 417728 99978 418048 100046
rect 417728 99922 417798 99978
rect 417854 99922 417922 99978
rect 417978 99922 418048 99978
rect 417728 99888 418048 99922
rect 420874 100350 421494 117922
rect 433088 112350 433408 112384
rect 433088 112294 433158 112350
rect 433214 112294 433282 112350
rect 433338 112294 433408 112350
rect 433088 112226 433408 112294
rect 433088 112170 433158 112226
rect 433214 112170 433282 112226
rect 433338 112170 433408 112226
rect 433088 112102 433408 112170
rect 433088 112046 433158 112102
rect 433214 112046 433282 112102
rect 433338 112046 433408 112102
rect 433088 111978 433408 112046
rect 433088 111922 433158 111978
rect 433214 111922 433282 111978
rect 433338 111922 433408 111978
rect 433088 111888 433408 111922
rect 435154 112350 435774 129922
rect 435154 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 435774 112350
rect 435154 112226 435774 112294
rect 435154 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 435774 112226
rect 435154 112102 435774 112170
rect 435154 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 435774 112102
rect 435154 111978 435774 112046
rect 435154 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 435774 111978
rect 420874 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 421494 100350
rect 420874 100226 421494 100294
rect 420874 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 421494 100226
rect 420874 100102 421494 100170
rect 420874 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 421494 100102
rect 420874 99978 421494 100046
rect 420874 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 421494 99978
rect 402874 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 403494 82350
rect 402874 82226 403494 82294
rect 402874 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 403494 82226
rect 402874 82102 403494 82170
rect 402874 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 403494 82102
rect 402874 81978 403494 82046
rect 402874 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 403494 81978
rect 399154 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 399774 76350
rect 399154 76226 399774 76294
rect 399154 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 399774 76226
rect 399154 76102 399774 76170
rect 399154 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 399774 76102
rect 399154 75978 399774 76046
rect 399154 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 399774 75978
rect 384874 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 385494 64350
rect 384874 64226 385494 64294
rect 384874 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 385494 64226
rect 384874 64102 385494 64170
rect 384874 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 385494 64102
rect 384874 63978 385494 64046
rect 384874 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 385494 63978
rect 384874 46350 385494 63922
rect 387008 64350 387328 64384
rect 387008 64294 387078 64350
rect 387134 64294 387202 64350
rect 387258 64294 387328 64350
rect 387008 64226 387328 64294
rect 387008 64170 387078 64226
rect 387134 64170 387202 64226
rect 387258 64170 387328 64226
rect 387008 64102 387328 64170
rect 387008 64046 387078 64102
rect 387134 64046 387202 64102
rect 387258 64046 387328 64102
rect 387008 63978 387328 64046
rect 387008 63922 387078 63978
rect 387134 63922 387202 63978
rect 387258 63922 387328 63978
rect 387008 63888 387328 63922
rect 384874 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 385494 46350
rect 384874 46226 385494 46294
rect 384874 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 385494 46226
rect 384874 46102 385494 46170
rect 384874 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 385494 46102
rect 384874 45978 385494 46046
rect 384874 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 385494 45978
rect 384874 28350 385494 45922
rect 384874 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 385494 28350
rect 384874 28226 385494 28294
rect 384874 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 385494 28226
rect 384874 28102 385494 28170
rect 384874 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 385494 28102
rect 384874 27978 385494 28046
rect 384874 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 385494 27978
rect 384874 10350 385494 27922
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 58350 399774 75922
rect 402368 76350 402688 76384
rect 402368 76294 402438 76350
rect 402494 76294 402562 76350
rect 402618 76294 402688 76350
rect 402368 76226 402688 76294
rect 402368 76170 402438 76226
rect 402494 76170 402562 76226
rect 402618 76170 402688 76226
rect 402368 76102 402688 76170
rect 402368 76046 402438 76102
rect 402494 76046 402562 76102
rect 402618 76046 402688 76102
rect 402368 75978 402688 76046
rect 402368 75922 402438 75978
rect 402494 75922 402562 75978
rect 402618 75922 402688 75978
rect 402368 75888 402688 75922
rect 399154 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 399774 58350
rect 399154 58226 399774 58294
rect 399154 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 399774 58226
rect 399154 58102 399774 58170
rect 399154 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 399774 58102
rect 399154 57978 399774 58046
rect 399154 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 399774 57978
rect 399154 40350 399774 57922
rect 399154 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 399774 40350
rect 399154 40226 399774 40294
rect 399154 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 399774 40226
rect 399154 40102 399774 40170
rect 399154 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 399774 40102
rect 399154 39978 399774 40046
rect 399154 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 399774 39978
rect 399154 22350 399774 39922
rect 399154 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 399774 22350
rect 399154 22226 399774 22294
rect 399154 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 399774 22226
rect 399154 22102 399774 22170
rect 399154 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 399774 22102
rect 399154 21978 399774 22046
rect 399154 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 399774 21978
rect 399154 4350 399774 21922
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 64350 403494 81922
rect 417728 82350 418048 82384
rect 417728 82294 417798 82350
rect 417854 82294 417922 82350
rect 417978 82294 418048 82350
rect 417728 82226 418048 82294
rect 417728 82170 417798 82226
rect 417854 82170 417922 82226
rect 417978 82170 418048 82226
rect 417728 82102 418048 82170
rect 417728 82046 417798 82102
rect 417854 82046 417922 82102
rect 417978 82046 418048 82102
rect 417728 81978 418048 82046
rect 417728 81922 417798 81978
rect 417854 81922 417922 81978
rect 417978 81922 418048 81978
rect 417728 81888 418048 81922
rect 420874 82350 421494 99922
rect 433088 94350 433408 94384
rect 433088 94294 433158 94350
rect 433214 94294 433282 94350
rect 433338 94294 433408 94350
rect 433088 94226 433408 94294
rect 433088 94170 433158 94226
rect 433214 94170 433282 94226
rect 433338 94170 433408 94226
rect 433088 94102 433408 94170
rect 433088 94046 433158 94102
rect 433214 94046 433282 94102
rect 433338 94046 433408 94102
rect 433088 93978 433408 94046
rect 433088 93922 433158 93978
rect 433214 93922 433282 93978
rect 433338 93922 433408 93978
rect 433088 93888 433408 93922
rect 435154 94350 435774 111922
rect 435154 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 435774 94350
rect 435154 94226 435774 94294
rect 435154 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 435774 94226
rect 435154 94102 435774 94170
rect 435154 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 435774 94102
rect 435154 93978 435774 94046
rect 435154 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 435774 93978
rect 420874 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 421494 82350
rect 420874 82226 421494 82294
rect 420874 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 421494 82226
rect 420874 82102 421494 82170
rect 420874 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 421494 82102
rect 420874 81978 421494 82046
rect 420874 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 421494 81978
rect 402874 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 403494 64350
rect 402874 64226 403494 64294
rect 402874 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 403494 64226
rect 402874 64102 403494 64170
rect 402874 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 403494 64102
rect 402874 63978 403494 64046
rect 402874 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 403494 63978
rect 402874 46350 403494 63922
rect 417728 64350 418048 64384
rect 417728 64294 417798 64350
rect 417854 64294 417922 64350
rect 417978 64294 418048 64350
rect 417728 64226 418048 64294
rect 417728 64170 417798 64226
rect 417854 64170 417922 64226
rect 417978 64170 418048 64226
rect 417728 64102 418048 64170
rect 417728 64046 417798 64102
rect 417854 64046 417922 64102
rect 417978 64046 418048 64102
rect 417728 63978 418048 64046
rect 417728 63922 417798 63978
rect 417854 63922 417922 63978
rect 417978 63922 418048 63978
rect 417728 63888 418048 63922
rect 420874 64350 421494 81922
rect 433088 76350 433408 76384
rect 433088 76294 433158 76350
rect 433214 76294 433282 76350
rect 433338 76294 433408 76350
rect 433088 76226 433408 76294
rect 433088 76170 433158 76226
rect 433214 76170 433282 76226
rect 433338 76170 433408 76226
rect 433088 76102 433408 76170
rect 433088 76046 433158 76102
rect 433214 76046 433282 76102
rect 433338 76046 433408 76102
rect 433088 75978 433408 76046
rect 433088 75922 433158 75978
rect 433214 75922 433282 75978
rect 433338 75922 433408 75978
rect 433088 75888 433408 75922
rect 435154 76350 435774 93922
rect 435154 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 435774 76350
rect 435154 76226 435774 76294
rect 435154 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 435774 76226
rect 435154 76102 435774 76170
rect 435154 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 435774 76102
rect 435154 75978 435774 76046
rect 435154 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 435774 75978
rect 420874 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 421494 64350
rect 420874 64226 421494 64294
rect 420874 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 421494 64226
rect 420874 64102 421494 64170
rect 420874 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 421494 64102
rect 420874 63978 421494 64046
rect 420874 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 421494 63978
rect 402874 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 403494 46350
rect 402874 46226 403494 46294
rect 402874 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 403494 46226
rect 402874 46102 403494 46170
rect 402874 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 403494 46102
rect 402874 45978 403494 46046
rect 402874 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 403494 45978
rect 402874 28350 403494 45922
rect 402874 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 403494 28350
rect 402874 28226 403494 28294
rect 402874 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 403494 28226
rect 402874 28102 403494 28170
rect 402874 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 403494 28102
rect 402874 27978 403494 28046
rect 402874 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 403494 27978
rect 402874 10350 403494 27922
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 58350 417774 61020
rect 417154 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 417774 58350
rect 417154 58226 417774 58294
rect 417154 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 417774 58226
rect 417154 58102 417774 58170
rect 417154 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 417774 58102
rect 417154 57978 417774 58046
rect 417154 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 417774 57978
rect 417154 40350 417774 57922
rect 417154 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 417774 40350
rect 417154 40226 417774 40294
rect 417154 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 417774 40226
rect 417154 40102 417774 40170
rect 417154 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 417774 40102
rect 417154 39978 417774 40046
rect 417154 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 417774 39978
rect 417154 22350 417774 39922
rect 417154 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 417774 22350
rect 417154 22226 417774 22294
rect 417154 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 417774 22226
rect 417154 22102 417774 22170
rect 417154 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 417774 22102
rect 417154 21978 417774 22046
rect 417154 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 417774 21978
rect 417154 4350 417774 21922
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 46350 421494 63922
rect 420874 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 421494 46350
rect 420874 46226 421494 46294
rect 420874 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 421494 46226
rect 420874 46102 421494 46170
rect 420874 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 421494 46102
rect 420874 45978 421494 46046
rect 420874 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 421494 45978
rect 420874 28350 421494 45922
rect 420874 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 421494 28350
rect 420874 28226 421494 28294
rect 420874 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 421494 28226
rect 420874 28102 421494 28170
rect 420874 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 421494 28102
rect 420874 27978 421494 28046
rect 420874 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 421494 27978
rect 420874 10350 421494 27922
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 58350 435774 75922
rect 435154 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 435774 58350
rect 435154 58226 435774 58294
rect 435154 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 435774 58226
rect 435154 58102 435774 58170
rect 435154 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 435774 58102
rect 435154 57978 435774 58046
rect 435154 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 435774 57978
rect 435154 40350 435774 57922
rect 435154 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 435774 40350
rect 435154 40226 435774 40294
rect 435154 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 435774 40226
rect 435154 40102 435774 40170
rect 435154 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 435774 40102
rect 435154 39978 435774 40046
rect 435154 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 435774 39978
rect 435154 22350 435774 39922
rect 435154 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 435774 22350
rect 435154 22226 435774 22294
rect 435154 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 435774 22226
rect 435154 22102 435774 22170
rect 435154 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 435774 22102
rect 435154 21978 435774 22046
rect 435154 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 435774 21978
rect 435154 4350 435774 21922
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 514350 439494 531922
rect 438874 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 439494 514350
rect 438874 514226 439494 514294
rect 438874 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 439494 514226
rect 438874 514102 439494 514170
rect 438874 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 439494 514102
rect 438874 513978 439494 514046
rect 438874 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 439494 513978
rect 438874 496350 439494 513922
rect 438874 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 439494 496350
rect 438874 496226 439494 496294
rect 438874 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 439494 496226
rect 438874 496102 439494 496170
rect 438874 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 439494 496102
rect 438874 495978 439494 496046
rect 438874 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 439494 495978
rect 438874 478350 439494 495922
rect 438874 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 439494 478350
rect 438874 478226 439494 478294
rect 438874 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 439494 478226
rect 438874 478102 439494 478170
rect 438874 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 439494 478102
rect 438874 477978 439494 478046
rect 438874 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 439494 477978
rect 438874 460350 439494 477922
rect 438874 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 439494 460350
rect 438874 460226 439494 460294
rect 438874 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 439494 460226
rect 438874 460102 439494 460170
rect 438874 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 439494 460102
rect 438874 459978 439494 460046
rect 438874 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 439494 459978
rect 438874 442350 439494 459922
rect 438874 442294 438970 442350
rect 439026 442294 439094 442350
rect 439150 442294 439218 442350
rect 439274 442294 439342 442350
rect 439398 442294 439494 442350
rect 438874 442226 439494 442294
rect 438874 442170 438970 442226
rect 439026 442170 439094 442226
rect 439150 442170 439218 442226
rect 439274 442170 439342 442226
rect 439398 442170 439494 442226
rect 438874 442102 439494 442170
rect 438874 442046 438970 442102
rect 439026 442046 439094 442102
rect 439150 442046 439218 442102
rect 439274 442046 439342 442102
rect 439398 442046 439494 442102
rect 438874 441978 439494 442046
rect 438874 441922 438970 441978
rect 439026 441922 439094 441978
rect 439150 441922 439218 441978
rect 439274 441922 439342 441978
rect 439398 441922 439494 441978
rect 438874 424350 439494 441922
rect 438874 424294 438970 424350
rect 439026 424294 439094 424350
rect 439150 424294 439218 424350
rect 439274 424294 439342 424350
rect 439398 424294 439494 424350
rect 438874 424226 439494 424294
rect 438874 424170 438970 424226
rect 439026 424170 439094 424226
rect 439150 424170 439218 424226
rect 439274 424170 439342 424226
rect 439398 424170 439494 424226
rect 438874 424102 439494 424170
rect 438874 424046 438970 424102
rect 439026 424046 439094 424102
rect 439150 424046 439218 424102
rect 439274 424046 439342 424102
rect 439398 424046 439494 424102
rect 438874 423978 439494 424046
rect 438874 423922 438970 423978
rect 439026 423922 439094 423978
rect 439150 423922 439218 423978
rect 439274 423922 439342 423978
rect 439398 423922 439494 423978
rect 438874 406350 439494 423922
rect 438874 406294 438970 406350
rect 439026 406294 439094 406350
rect 439150 406294 439218 406350
rect 439274 406294 439342 406350
rect 439398 406294 439494 406350
rect 438874 406226 439494 406294
rect 438874 406170 438970 406226
rect 439026 406170 439094 406226
rect 439150 406170 439218 406226
rect 439274 406170 439342 406226
rect 439398 406170 439494 406226
rect 438874 406102 439494 406170
rect 438874 406046 438970 406102
rect 439026 406046 439094 406102
rect 439150 406046 439218 406102
rect 439274 406046 439342 406102
rect 439398 406046 439494 406102
rect 438874 405978 439494 406046
rect 438874 405922 438970 405978
rect 439026 405922 439094 405978
rect 439150 405922 439218 405978
rect 439274 405922 439342 405978
rect 439398 405922 439494 405978
rect 438874 388350 439494 405922
rect 438874 388294 438970 388350
rect 439026 388294 439094 388350
rect 439150 388294 439218 388350
rect 439274 388294 439342 388350
rect 439398 388294 439494 388350
rect 438874 388226 439494 388294
rect 438874 388170 438970 388226
rect 439026 388170 439094 388226
rect 439150 388170 439218 388226
rect 439274 388170 439342 388226
rect 439398 388170 439494 388226
rect 438874 388102 439494 388170
rect 438874 388046 438970 388102
rect 439026 388046 439094 388102
rect 439150 388046 439218 388102
rect 439274 388046 439342 388102
rect 439398 388046 439494 388102
rect 438874 387978 439494 388046
rect 438874 387922 438970 387978
rect 439026 387922 439094 387978
rect 439150 387922 439218 387978
rect 439274 387922 439342 387978
rect 439398 387922 439494 387978
rect 438874 370350 439494 387922
rect 438874 370294 438970 370350
rect 439026 370294 439094 370350
rect 439150 370294 439218 370350
rect 439274 370294 439342 370350
rect 439398 370294 439494 370350
rect 438874 370226 439494 370294
rect 438874 370170 438970 370226
rect 439026 370170 439094 370226
rect 439150 370170 439218 370226
rect 439274 370170 439342 370226
rect 439398 370170 439494 370226
rect 438874 370102 439494 370170
rect 438874 370046 438970 370102
rect 439026 370046 439094 370102
rect 439150 370046 439218 370102
rect 439274 370046 439342 370102
rect 439398 370046 439494 370102
rect 438874 369978 439494 370046
rect 438874 369922 438970 369978
rect 439026 369922 439094 369978
rect 439150 369922 439218 369978
rect 439274 369922 439342 369978
rect 439398 369922 439494 369978
rect 438874 352350 439494 369922
rect 438874 352294 438970 352350
rect 439026 352294 439094 352350
rect 439150 352294 439218 352350
rect 439274 352294 439342 352350
rect 439398 352294 439494 352350
rect 438874 352226 439494 352294
rect 438874 352170 438970 352226
rect 439026 352170 439094 352226
rect 439150 352170 439218 352226
rect 439274 352170 439342 352226
rect 439398 352170 439494 352226
rect 438874 352102 439494 352170
rect 438874 352046 438970 352102
rect 439026 352046 439094 352102
rect 439150 352046 439218 352102
rect 439274 352046 439342 352102
rect 439398 352046 439494 352102
rect 438874 351978 439494 352046
rect 438874 351922 438970 351978
rect 439026 351922 439094 351978
rect 439150 351922 439218 351978
rect 439274 351922 439342 351978
rect 439398 351922 439494 351978
rect 438874 334350 439494 351922
rect 438874 334294 438970 334350
rect 439026 334294 439094 334350
rect 439150 334294 439218 334350
rect 439274 334294 439342 334350
rect 439398 334294 439494 334350
rect 438874 334226 439494 334294
rect 438874 334170 438970 334226
rect 439026 334170 439094 334226
rect 439150 334170 439218 334226
rect 439274 334170 439342 334226
rect 439398 334170 439494 334226
rect 438874 334102 439494 334170
rect 438874 334046 438970 334102
rect 439026 334046 439094 334102
rect 439150 334046 439218 334102
rect 439274 334046 439342 334102
rect 439398 334046 439494 334102
rect 438874 333978 439494 334046
rect 438874 333922 438970 333978
rect 439026 333922 439094 333978
rect 439150 333922 439218 333978
rect 439274 333922 439342 333978
rect 439398 333922 439494 333978
rect 438874 316350 439494 333922
rect 438874 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 439494 316350
rect 438874 316226 439494 316294
rect 438874 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 439494 316226
rect 438874 316102 439494 316170
rect 438874 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 439494 316102
rect 438874 315978 439494 316046
rect 438874 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 439494 315978
rect 438874 298350 439494 315922
rect 438874 298294 438970 298350
rect 439026 298294 439094 298350
rect 439150 298294 439218 298350
rect 439274 298294 439342 298350
rect 439398 298294 439494 298350
rect 438874 298226 439494 298294
rect 438874 298170 438970 298226
rect 439026 298170 439094 298226
rect 439150 298170 439218 298226
rect 439274 298170 439342 298226
rect 439398 298170 439494 298226
rect 438874 298102 439494 298170
rect 438874 298046 438970 298102
rect 439026 298046 439094 298102
rect 439150 298046 439218 298102
rect 439274 298046 439342 298102
rect 439398 298046 439494 298102
rect 438874 297978 439494 298046
rect 438874 297922 438970 297978
rect 439026 297922 439094 297978
rect 439150 297922 439218 297978
rect 439274 297922 439342 297978
rect 439398 297922 439494 297978
rect 438874 280350 439494 297922
rect 438874 280294 438970 280350
rect 439026 280294 439094 280350
rect 439150 280294 439218 280350
rect 439274 280294 439342 280350
rect 439398 280294 439494 280350
rect 438874 280226 439494 280294
rect 438874 280170 438970 280226
rect 439026 280170 439094 280226
rect 439150 280170 439218 280226
rect 439274 280170 439342 280226
rect 439398 280170 439494 280226
rect 438874 280102 439494 280170
rect 438874 280046 438970 280102
rect 439026 280046 439094 280102
rect 439150 280046 439218 280102
rect 439274 280046 439342 280102
rect 439398 280046 439494 280102
rect 438874 279978 439494 280046
rect 438874 279922 438970 279978
rect 439026 279922 439094 279978
rect 439150 279922 439218 279978
rect 439274 279922 439342 279978
rect 439398 279922 439494 279978
rect 438874 262350 439494 279922
rect 438874 262294 438970 262350
rect 439026 262294 439094 262350
rect 439150 262294 439218 262350
rect 439274 262294 439342 262350
rect 439398 262294 439494 262350
rect 438874 262226 439494 262294
rect 438874 262170 438970 262226
rect 439026 262170 439094 262226
rect 439150 262170 439218 262226
rect 439274 262170 439342 262226
rect 439398 262170 439494 262226
rect 438874 262102 439494 262170
rect 438874 262046 438970 262102
rect 439026 262046 439094 262102
rect 439150 262046 439218 262102
rect 439274 262046 439342 262102
rect 439398 262046 439494 262102
rect 438874 261978 439494 262046
rect 438874 261922 438970 261978
rect 439026 261922 439094 261978
rect 439150 261922 439218 261978
rect 439274 261922 439342 261978
rect 439398 261922 439494 261978
rect 438874 244350 439494 261922
rect 438874 244294 438970 244350
rect 439026 244294 439094 244350
rect 439150 244294 439218 244350
rect 439274 244294 439342 244350
rect 439398 244294 439494 244350
rect 438874 244226 439494 244294
rect 438874 244170 438970 244226
rect 439026 244170 439094 244226
rect 439150 244170 439218 244226
rect 439274 244170 439342 244226
rect 439398 244170 439494 244226
rect 438874 244102 439494 244170
rect 438874 244046 438970 244102
rect 439026 244046 439094 244102
rect 439150 244046 439218 244102
rect 439274 244046 439342 244102
rect 439398 244046 439494 244102
rect 438874 243978 439494 244046
rect 438874 243922 438970 243978
rect 439026 243922 439094 243978
rect 439150 243922 439218 243978
rect 439274 243922 439342 243978
rect 439398 243922 439494 243978
rect 438874 226350 439494 243922
rect 438874 226294 438970 226350
rect 439026 226294 439094 226350
rect 439150 226294 439218 226350
rect 439274 226294 439342 226350
rect 439398 226294 439494 226350
rect 438874 226226 439494 226294
rect 438874 226170 438970 226226
rect 439026 226170 439094 226226
rect 439150 226170 439218 226226
rect 439274 226170 439342 226226
rect 439398 226170 439494 226226
rect 438874 226102 439494 226170
rect 438874 226046 438970 226102
rect 439026 226046 439094 226102
rect 439150 226046 439218 226102
rect 439274 226046 439342 226102
rect 439398 226046 439494 226102
rect 438874 225978 439494 226046
rect 438874 225922 438970 225978
rect 439026 225922 439094 225978
rect 439150 225922 439218 225978
rect 439274 225922 439342 225978
rect 439398 225922 439494 225978
rect 438874 208350 439494 225922
rect 438874 208294 438970 208350
rect 439026 208294 439094 208350
rect 439150 208294 439218 208350
rect 439274 208294 439342 208350
rect 439398 208294 439494 208350
rect 438874 208226 439494 208294
rect 438874 208170 438970 208226
rect 439026 208170 439094 208226
rect 439150 208170 439218 208226
rect 439274 208170 439342 208226
rect 439398 208170 439494 208226
rect 438874 208102 439494 208170
rect 438874 208046 438970 208102
rect 439026 208046 439094 208102
rect 439150 208046 439218 208102
rect 439274 208046 439342 208102
rect 439398 208046 439494 208102
rect 438874 207978 439494 208046
rect 438874 207922 438970 207978
rect 439026 207922 439094 207978
rect 439150 207922 439218 207978
rect 439274 207922 439342 207978
rect 439398 207922 439494 207978
rect 438874 190350 439494 207922
rect 438874 190294 438970 190350
rect 439026 190294 439094 190350
rect 439150 190294 439218 190350
rect 439274 190294 439342 190350
rect 439398 190294 439494 190350
rect 438874 190226 439494 190294
rect 438874 190170 438970 190226
rect 439026 190170 439094 190226
rect 439150 190170 439218 190226
rect 439274 190170 439342 190226
rect 439398 190170 439494 190226
rect 438874 190102 439494 190170
rect 438874 190046 438970 190102
rect 439026 190046 439094 190102
rect 439150 190046 439218 190102
rect 439274 190046 439342 190102
rect 439398 190046 439494 190102
rect 438874 189978 439494 190046
rect 438874 189922 438970 189978
rect 439026 189922 439094 189978
rect 439150 189922 439218 189978
rect 439274 189922 439342 189978
rect 439398 189922 439494 189978
rect 438874 172350 439494 189922
rect 438874 172294 438970 172350
rect 439026 172294 439094 172350
rect 439150 172294 439218 172350
rect 439274 172294 439342 172350
rect 439398 172294 439494 172350
rect 438874 172226 439494 172294
rect 438874 172170 438970 172226
rect 439026 172170 439094 172226
rect 439150 172170 439218 172226
rect 439274 172170 439342 172226
rect 439398 172170 439494 172226
rect 438874 172102 439494 172170
rect 438874 172046 438970 172102
rect 439026 172046 439094 172102
rect 439150 172046 439218 172102
rect 439274 172046 439342 172102
rect 439398 172046 439494 172102
rect 438874 171978 439494 172046
rect 438874 171922 438970 171978
rect 439026 171922 439094 171978
rect 439150 171922 439218 171978
rect 439274 171922 439342 171978
rect 439398 171922 439494 171978
rect 438874 154350 439494 171922
rect 438874 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 439494 154350
rect 438874 154226 439494 154294
rect 438874 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 439494 154226
rect 438874 154102 439494 154170
rect 438874 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 439494 154102
rect 438874 153978 439494 154046
rect 438874 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 439494 153978
rect 438874 136350 439494 153922
rect 438874 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 439494 136350
rect 438874 136226 439494 136294
rect 438874 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 439494 136226
rect 438874 136102 439494 136170
rect 438874 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 439494 136102
rect 438874 135978 439494 136046
rect 438874 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 439494 135978
rect 438874 118350 439494 135922
rect 438874 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 439494 118350
rect 438874 118226 439494 118294
rect 438874 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 439494 118226
rect 438874 118102 439494 118170
rect 438874 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 439494 118102
rect 438874 117978 439494 118046
rect 438874 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 439494 117978
rect 438874 100350 439494 117922
rect 438874 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 439494 100350
rect 438874 100226 439494 100294
rect 438874 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 439494 100226
rect 438874 100102 439494 100170
rect 438874 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 439494 100102
rect 438874 99978 439494 100046
rect 438874 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 439494 99978
rect 438874 82350 439494 99922
rect 438874 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 439494 82350
rect 438874 82226 439494 82294
rect 438874 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 439494 82226
rect 438874 82102 439494 82170
rect 438874 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 439494 82102
rect 438874 81978 439494 82046
rect 438874 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 439494 81978
rect 438874 64350 439494 81922
rect 438874 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 439494 64350
rect 438874 64226 439494 64294
rect 438874 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 439494 64226
rect 438874 64102 439494 64170
rect 438874 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 439494 64102
rect 438874 63978 439494 64046
rect 438874 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 439494 63978
rect 438874 46350 439494 63922
rect 438874 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 439494 46350
rect 438874 46226 439494 46294
rect 438874 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 439494 46226
rect 438874 46102 439494 46170
rect 438874 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 439494 46102
rect 438874 45978 439494 46046
rect 438874 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 439494 45978
rect 438874 28350 439494 45922
rect 438874 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 439494 28350
rect 438874 28226 439494 28294
rect 438874 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 439494 28226
rect 438874 28102 439494 28170
rect 438874 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 439494 28102
rect 438874 27978 439494 28046
rect 438874 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 439494 27978
rect 438874 10350 439494 27922
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 526350 453774 543922
rect 453154 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 453774 526350
rect 453154 526226 453774 526294
rect 453154 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 453774 526226
rect 453154 526102 453774 526170
rect 453154 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 453774 526102
rect 453154 525978 453774 526046
rect 453154 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 453774 525978
rect 453154 508350 453774 525922
rect 453154 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 453774 508350
rect 453154 508226 453774 508294
rect 453154 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 453774 508226
rect 453154 508102 453774 508170
rect 453154 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 453774 508102
rect 453154 507978 453774 508046
rect 453154 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 453774 507978
rect 453154 490350 453774 507922
rect 453154 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 453774 490350
rect 453154 490226 453774 490294
rect 453154 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 453774 490226
rect 453154 490102 453774 490170
rect 453154 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 453774 490102
rect 453154 489978 453774 490046
rect 453154 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 453774 489978
rect 453154 472350 453774 489922
rect 453154 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 453774 472350
rect 453154 472226 453774 472294
rect 453154 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 453774 472226
rect 453154 472102 453774 472170
rect 453154 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 453774 472102
rect 453154 471978 453774 472046
rect 453154 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 453774 471978
rect 453154 454350 453774 471922
rect 453154 454294 453250 454350
rect 453306 454294 453374 454350
rect 453430 454294 453498 454350
rect 453554 454294 453622 454350
rect 453678 454294 453774 454350
rect 453154 454226 453774 454294
rect 453154 454170 453250 454226
rect 453306 454170 453374 454226
rect 453430 454170 453498 454226
rect 453554 454170 453622 454226
rect 453678 454170 453774 454226
rect 453154 454102 453774 454170
rect 453154 454046 453250 454102
rect 453306 454046 453374 454102
rect 453430 454046 453498 454102
rect 453554 454046 453622 454102
rect 453678 454046 453774 454102
rect 453154 453978 453774 454046
rect 453154 453922 453250 453978
rect 453306 453922 453374 453978
rect 453430 453922 453498 453978
rect 453554 453922 453622 453978
rect 453678 453922 453774 453978
rect 453154 436350 453774 453922
rect 453154 436294 453250 436350
rect 453306 436294 453374 436350
rect 453430 436294 453498 436350
rect 453554 436294 453622 436350
rect 453678 436294 453774 436350
rect 453154 436226 453774 436294
rect 453154 436170 453250 436226
rect 453306 436170 453374 436226
rect 453430 436170 453498 436226
rect 453554 436170 453622 436226
rect 453678 436170 453774 436226
rect 453154 436102 453774 436170
rect 453154 436046 453250 436102
rect 453306 436046 453374 436102
rect 453430 436046 453498 436102
rect 453554 436046 453622 436102
rect 453678 436046 453774 436102
rect 453154 435978 453774 436046
rect 453154 435922 453250 435978
rect 453306 435922 453374 435978
rect 453430 435922 453498 435978
rect 453554 435922 453622 435978
rect 453678 435922 453774 435978
rect 453154 418350 453774 435922
rect 453154 418294 453250 418350
rect 453306 418294 453374 418350
rect 453430 418294 453498 418350
rect 453554 418294 453622 418350
rect 453678 418294 453774 418350
rect 453154 418226 453774 418294
rect 453154 418170 453250 418226
rect 453306 418170 453374 418226
rect 453430 418170 453498 418226
rect 453554 418170 453622 418226
rect 453678 418170 453774 418226
rect 453154 418102 453774 418170
rect 453154 418046 453250 418102
rect 453306 418046 453374 418102
rect 453430 418046 453498 418102
rect 453554 418046 453622 418102
rect 453678 418046 453774 418102
rect 453154 417978 453774 418046
rect 453154 417922 453250 417978
rect 453306 417922 453374 417978
rect 453430 417922 453498 417978
rect 453554 417922 453622 417978
rect 453678 417922 453774 417978
rect 453154 400350 453774 417922
rect 453154 400294 453250 400350
rect 453306 400294 453374 400350
rect 453430 400294 453498 400350
rect 453554 400294 453622 400350
rect 453678 400294 453774 400350
rect 453154 400226 453774 400294
rect 453154 400170 453250 400226
rect 453306 400170 453374 400226
rect 453430 400170 453498 400226
rect 453554 400170 453622 400226
rect 453678 400170 453774 400226
rect 453154 400102 453774 400170
rect 453154 400046 453250 400102
rect 453306 400046 453374 400102
rect 453430 400046 453498 400102
rect 453554 400046 453622 400102
rect 453678 400046 453774 400102
rect 453154 399978 453774 400046
rect 453154 399922 453250 399978
rect 453306 399922 453374 399978
rect 453430 399922 453498 399978
rect 453554 399922 453622 399978
rect 453678 399922 453774 399978
rect 453154 382350 453774 399922
rect 453154 382294 453250 382350
rect 453306 382294 453374 382350
rect 453430 382294 453498 382350
rect 453554 382294 453622 382350
rect 453678 382294 453774 382350
rect 453154 382226 453774 382294
rect 453154 382170 453250 382226
rect 453306 382170 453374 382226
rect 453430 382170 453498 382226
rect 453554 382170 453622 382226
rect 453678 382170 453774 382226
rect 453154 382102 453774 382170
rect 453154 382046 453250 382102
rect 453306 382046 453374 382102
rect 453430 382046 453498 382102
rect 453554 382046 453622 382102
rect 453678 382046 453774 382102
rect 453154 381978 453774 382046
rect 453154 381922 453250 381978
rect 453306 381922 453374 381978
rect 453430 381922 453498 381978
rect 453554 381922 453622 381978
rect 453678 381922 453774 381978
rect 453154 364350 453774 381922
rect 453154 364294 453250 364350
rect 453306 364294 453374 364350
rect 453430 364294 453498 364350
rect 453554 364294 453622 364350
rect 453678 364294 453774 364350
rect 453154 364226 453774 364294
rect 453154 364170 453250 364226
rect 453306 364170 453374 364226
rect 453430 364170 453498 364226
rect 453554 364170 453622 364226
rect 453678 364170 453774 364226
rect 453154 364102 453774 364170
rect 453154 364046 453250 364102
rect 453306 364046 453374 364102
rect 453430 364046 453498 364102
rect 453554 364046 453622 364102
rect 453678 364046 453774 364102
rect 453154 363978 453774 364046
rect 453154 363922 453250 363978
rect 453306 363922 453374 363978
rect 453430 363922 453498 363978
rect 453554 363922 453622 363978
rect 453678 363922 453774 363978
rect 453154 346350 453774 363922
rect 453154 346294 453250 346350
rect 453306 346294 453374 346350
rect 453430 346294 453498 346350
rect 453554 346294 453622 346350
rect 453678 346294 453774 346350
rect 453154 346226 453774 346294
rect 453154 346170 453250 346226
rect 453306 346170 453374 346226
rect 453430 346170 453498 346226
rect 453554 346170 453622 346226
rect 453678 346170 453774 346226
rect 453154 346102 453774 346170
rect 453154 346046 453250 346102
rect 453306 346046 453374 346102
rect 453430 346046 453498 346102
rect 453554 346046 453622 346102
rect 453678 346046 453774 346102
rect 453154 345978 453774 346046
rect 453154 345922 453250 345978
rect 453306 345922 453374 345978
rect 453430 345922 453498 345978
rect 453554 345922 453622 345978
rect 453678 345922 453774 345978
rect 453154 328350 453774 345922
rect 453154 328294 453250 328350
rect 453306 328294 453374 328350
rect 453430 328294 453498 328350
rect 453554 328294 453622 328350
rect 453678 328294 453774 328350
rect 453154 328226 453774 328294
rect 453154 328170 453250 328226
rect 453306 328170 453374 328226
rect 453430 328170 453498 328226
rect 453554 328170 453622 328226
rect 453678 328170 453774 328226
rect 453154 328102 453774 328170
rect 453154 328046 453250 328102
rect 453306 328046 453374 328102
rect 453430 328046 453498 328102
rect 453554 328046 453622 328102
rect 453678 328046 453774 328102
rect 453154 327978 453774 328046
rect 453154 327922 453250 327978
rect 453306 327922 453374 327978
rect 453430 327922 453498 327978
rect 453554 327922 453622 327978
rect 453678 327922 453774 327978
rect 453154 310350 453774 327922
rect 453154 310294 453250 310350
rect 453306 310294 453374 310350
rect 453430 310294 453498 310350
rect 453554 310294 453622 310350
rect 453678 310294 453774 310350
rect 453154 310226 453774 310294
rect 453154 310170 453250 310226
rect 453306 310170 453374 310226
rect 453430 310170 453498 310226
rect 453554 310170 453622 310226
rect 453678 310170 453774 310226
rect 453154 310102 453774 310170
rect 453154 310046 453250 310102
rect 453306 310046 453374 310102
rect 453430 310046 453498 310102
rect 453554 310046 453622 310102
rect 453678 310046 453774 310102
rect 453154 309978 453774 310046
rect 453154 309922 453250 309978
rect 453306 309922 453374 309978
rect 453430 309922 453498 309978
rect 453554 309922 453622 309978
rect 453678 309922 453774 309978
rect 453154 292350 453774 309922
rect 453154 292294 453250 292350
rect 453306 292294 453374 292350
rect 453430 292294 453498 292350
rect 453554 292294 453622 292350
rect 453678 292294 453774 292350
rect 453154 292226 453774 292294
rect 453154 292170 453250 292226
rect 453306 292170 453374 292226
rect 453430 292170 453498 292226
rect 453554 292170 453622 292226
rect 453678 292170 453774 292226
rect 453154 292102 453774 292170
rect 453154 292046 453250 292102
rect 453306 292046 453374 292102
rect 453430 292046 453498 292102
rect 453554 292046 453622 292102
rect 453678 292046 453774 292102
rect 453154 291978 453774 292046
rect 453154 291922 453250 291978
rect 453306 291922 453374 291978
rect 453430 291922 453498 291978
rect 453554 291922 453622 291978
rect 453678 291922 453774 291978
rect 453154 274350 453774 291922
rect 453154 274294 453250 274350
rect 453306 274294 453374 274350
rect 453430 274294 453498 274350
rect 453554 274294 453622 274350
rect 453678 274294 453774 274350
rect 453154 274226 453774 274294
rect 453154 274170 453250 274226
rect 453306 274170 453374 274226
rect 453430 274170 453498 274226
rect 453554 274170 453622 274226
rect 453678 274170 453774 274226
rect 453154 274102 453774 274170
rect 453154 274046 453250 274102
rect 453306 274046 453374 274102
rect 453430 274046 453498 274102
rect 453554 274046 453622 274102
rect 453678 274046 453774 274102
rect 453154 273978 453774 274046
rect 453154 273922 453250 273978
rect 453306 273922 453374 273978
rect 453430 273922 453498 273978
rect 453554 273922 453622 273978
rect 453678 273922 453774 273978
rect 453154 256350 453774 273922
rect 453154 256294 453250 256350
rect 453306 256294 453374 256350
rect 453430 256294 453498 256350
rect 453554 256294 453622 256350
rect 453678 256294 453774 256350
rect 453154 256226 453774 256294
rect 453154 256170 453250 256226
rect 453306 256170 453374 256226
rect 453430 256170 453498 256226
rect 453554 256170 453622 256226
rect 453678 256170 453774 256226
rect 453154 256102 453774 256170
rect 453154 256046 453250 256102
rect 453306 256046 453374 256102
rect 453430 256046 453498 256102
rect 453554 256046 453622 256102
rect 453678 256046 453774 256102
rect 453154 255978 453774 256046
rect 453154 255922 453250 255978
rect 453306 255922 453374 255978
rect 453430 255922 453498 255978
rect 453554 255922 453622 255978
rect 453678 255922 453774 255978
rect 453154 238350 453774 255922
rect 453154 238294 453250 238350
rect 453306 238294 453374 238350
rect 453430 238294 453498 238350
rect 453554 238294 453622 238350
rect 453678 238294 453774 238350
rect 453154 238226 453774 238294
rect 453154 238170 453250 238226
rect 453306 238170 453374 238226
rect 453430 238170 453498 238226
rect 453554 238170 453622 238226
rect 453678 238170 453774 238226
rect 453154 238102 453774 238170
rect 453154 238046 453250 238102
rect 453306 238046 453374 238102
rect 453430 238046 453498 238102
rect 453554 238046 453622 238102
rect 453678 238046 453774 238102
rect 453154 237978 453774 238046
rect 453154 237922 453250 237978
rect 453306 237922 453374 237978
rect 453430 237922 453498 237978
rect 453554 237922 453622 237978
rect 453678 237922 453774 237978
rect 453154 220350 453774 237922
rect 453154 220294 453250 220350
rect 453306 220294 453374 220350
rect 453430 220294 453498 220350
rect 453554 220294 453622 220350
rect 453678 220294 453774 220350
rect 453154 220226 453774 220294
rect 453154 220170 453250 220226
rect 453306 220170 453374 220226
rect 453430 220170 453498 220226
rect 453554 220170 453622 220226
rect 453678 220170 453774 220226
rect 453154 220102 453774 220170
rect 453154 220046 453250 220102
rect 453306 220046 453374 220102
rect 453430 220046 453498 220102
rect 453554 220046 453622 220102
rect 453678 220046 453774 220102
rect 453154 219978 453774 220046
rect 453154 219922 453250 219978
rect 453306 219922 453374 219978
rect 453430 219922 453498 219978
rect 453554 219922 453622 219978
rect 453678 219922 453774 219978
rect 453154 202350 453774 219922
rect 453154 202294 453250 202350
rect 453306 202294 453374 202350
rect 453430 202294 453498 202350
rect 453554 202294 453622 202350
rect 453678 202294 453774 202350
rect 453154 202226 453774 202294
rect 453154 202170 453250 202226
rect 453306 202170 453374 202226
rect 453430 202170 453498 202226
rect 453554 202170 453622 202226
rect 453678 202170 453774 202226
rect 453154 202102 453774 202170
rect 453154 202046 453250 202102
rect 453306 202046 453374 202102
rect 453430 202046 453498 202102
rect 453554 202046 453622 202102
rect 453678 202046 453774 202102
rect 453154 201978 453774 202046
rect 453154 201922 453250 201978
rect 453306 201922 453374 201978
rect 453430 201922 453498 201978
rect 453554 201922 453622 201978
rect 453678 201922 453774 201978
rect 453154 184350 453774 201922
rect 453154 184294 453250 184350
rect 453306 184294 453374 184350
rect 453430 184294 453498 184350
rect 453554 184294 453622 184350
rect 453678 184294 453774 184350
rect 453154 184226 453774 184294
rect 453154 184170 453250 184226
rect 453306 184170 453374 184226
rect 453430 184170 453498 184226
rect 453554 184170 453622 184226
rect 453678 184170 453774 184226
rect 453154 184102 453774 184170
rect 453154 184046 453250 184102
rect 453306 184046 453374 184102
rect 453430 184046 453498 184102
rect 453554 184046 453622 184102
rect 453678 184046 453774 184102
rect 453154 183978 453774 184046
rect 453154 183922 453250 183978
rect 453306 183922 453374 183978
rect 453430 183922 453498 183978
rect 453554 183922 453622 183978
rect 453678 183922 453774 183978
rect 453154 166350 453774 183922
rect 453154 166294 453250 166350
rect 453306 166294 453374 166350
rect 453430 166294 453498 166350
rect 453554 166294 453622 166350
rect 453678 166294 453774 166350
rect 453154 166226 453774 166294
rect 453154 166170 453250 166226
rect 453306 166170 453374 166226
rect 453430 166170 453498 166226
rect 453554 166170 453622 166226
rect 453678 166170 453774 166226
rect 453154 166102 453774 166170
rect 453154 166046 453250 166102
rect 453306 166046 453374 166102
rect 453430 166046 453498 166102
rect 453554 166046 453622 166102
rect 453678 166046 453774 166102
rect 453154 165978 453774 166046
rect 453154 165922 453250 165978
rect 453306 165922 453374 165978
rect 453430 165922 453498 165978
rect 453554 165922 453622 165978
rect 453678 165922 453774 165978
rect 453154 148350 453774 165922
rect 453154 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 453774 148350
rect 453154 148226 453774 148294
rect 453154 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 453774 148226
rect 453154 148102 453774 148170
rect 453154 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 453774 148102
rect 453154 147978 453774 148046
rect 453154 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 453774 147978
rect 453154 130350 453774 147922
rect 453154 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 453774 130350
rect 453154 130226 453774 130294
rect 453154 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 453774 130226
rect 453154 130102 453774 130170
rect 453154 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 453774 130102
rect 453154 129978 453774 130046
rect 453154 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 453774 129978
rect 453154 112350 453774 129922
rect 453154 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 453774 112350
rect 453154 112226 453774 112294
rect 453154 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 453774 112226
rect 453154 112102 453774 112170
rect 453154 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 453774 112102
rect 453154 111978 453774 112046
rect 453154 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 453774 111978
rect 453154 94350 453774 111922
rect 453154 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 453774 94350
rect 453154 94226 453774 94294
rect 453154 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 453774 94226
rect 453154 94102 453774 94170
rect 453154 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 453774 94102
rect 453154 93978 453774 94046
rect 453154 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 453774 93978
rect 453154 76350 453774 93922
rect 453154 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 453774 76350
rect 453154 76226 453774 76294
rect 453154 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 453774 76226
rect 453154 76102 453774 76170
rect 453154 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 453774 76102
rect 453154 75978 453774 76046
rect 453154 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 453774 75978
rect 453154 58350 453774 75922
rect 453154 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 453774 58350
rect 453154 58226 453774 58294
rect 453154 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 453774 58226
rect 453154 58102 453774 58170
rect 453154 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 453774 58102
rect 453154 57978 453774 58046
rect 453154 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 453774 57978
rect 453154 40350 453774 57922
rect 453154 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 453774 40350
rect 453154 40226 453774 40294
rect 453154 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 453774 40226
rect 453154 40102 453774 40170
rect 453154 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 453774 40102
rect 453154 39978 453774 40046
rect 453154 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 453774 39978
rect 453154 22350 453774 39922
rect 453154 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 453774 22350
rect 453154 22226 453774 22294
rect 453154 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 453774 22226
rect 453154 22102 453774 22170
rect 453154 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 453774 22102
rect 453154 21978 453774 22046
rect 453154 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 453774 21978
rect 453154 4350 453774 21922
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 514350 457494 531922
rect 456874 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 457494 514350
rect 456874 514226 457494 514294
rect 456874 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 457494 514226
rect 456874 514102 457494 514170
rect 456874 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 457494 514102
rect 456874 513978 457494 514046
rect 456874 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 457494 513978
rect 456874 496350 457494 513922
rect 456874 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 457494 496350
rect 456874 496226 457494 496294
rect 456874 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 457494 496226
rect 456874 496102 457494 496170
rect 456874 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 457494 496102
rect 456874 495978 457494 496046
rect 456874 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 457494 495978
rect 456874 478350 457494 495922
rect 456874 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 457494 478350
rect 456874 478226 457494 478294
rect 456874 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 457494 478226
rect 456874 478102 457494 478170
rect 456874 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 457494 478102
rect 456874 477978 457494 478046
rect 456874 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 457494 477978
rect 456874 460350 457494 477922
rect 456874 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 457494 460350
rect 456874 460226 457494 460294
rect 456874 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 457494 460226
rect 456874 460102 457494 460170
rect 456874 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 457494 460102
rect 456874 459978 457494 460046
rect 456874 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 457494 459978
rect 456874 442350 457494 459922
rect 456874 442294 456970 442350
rect 457026 442294 457094 442350
rect 457150 442294 457218 442350
rect 457274 442294 457342 442350
rect 457398 442294 457494 442350
rect 456874 442226 457494 442294
rect 456874 442170 456970 442226
rect 457026 442170 457094 442226
rect 457150 442170 457218 442226
rect 457274 442170 457342 442226
rect 457398 442170 457494 442226
rect 456874 442102 457494 442170
rect 456874 442046 456970 442102
rect 457026 442046 457094 442102
rect 457150 442046 457218 442102
rect 457274 442046 457342 442102
rect 457398 442046 457494 442102
rect 456874 441978 457494 442046
rect 456874 441922 456970 441978
rect 457026 441922 457094 441978
rect 457150 441922 457218 441978
rect 457274 441922 457342 441978
rect 457398 441922 457494 441978
rect 456874 424350 457494 441922
rect 456874 424294 456970 424350
rect 457026 424294 457094 424350
rect 457150 424294 457218 424350
rect 457274 424294 457342 424350
rect 457398 424294 457494 424350
rect 456874 424226 457494 424294
rect 456874 424170 456970 424226
rect 457026 424170 457094 424226
rect 457150 424170 457218 424226
rect 457274 424170 457342 424226
rect 457398 424170 457494 424226
rect 456874 424102 457494 424170
rect 456874 424046 456970 424102
rect 457026 424046 457094 424102
rect 457150 424046 457218 424102
rect 457274 424046 457342 424102
rect 457398 424046 457494 424102
rect 456874 423978 457494 424046
rect 456874 423922 456970 423978
rect 457026 423922 457094 423978
rect 457150 423922 457218 423978
rect 457274 423922 457342 423978
rect 457398 423922 457494 423978
rect 456874 406350 457494 423922
rect 456874 406294 456970 406350
rect 457026 406294 457094 406350
rect 457150 406294 457218 406350
rect 457274 406294 457342 406350
rect 457398 406294 457494 406350
rect 456874 406226 457494 406294
rect 456874 406170 456970 406226
rect 457026 406170 457094 406226
rect 457150 406170 457218 406226
rect 457274 406170 457342 406226
rect 457398 406170 457494 406226
rect 456874 406102 457494 406170
rect 456874 406046 456970 406102
rect 457026 406046 457094 406102
rect 457150 406046 457218 406102
rect 457274 406046 457342 406102
rect 457398 406046 457494 406102
rect 456874 405978 457494 406046
rect 456874 405922 456970 405978
rect 457026 405922 457094 405978
rect 457150 405922 457218 405978
rect 457274 405922 457342 405978
rect 457398 405922 457494 405978
rect 456874 388350 457494 405922
rect 456874 388294 456970 388350
rect 457026 388294 457094 388350
rect 457150 388294 457218 388350
rect 457274 388294 457342 388350
rect 457398 388294 457494 388350
rect 456874 388226 457494 388294
rect 456874 388170 456970 388226
rect 457026 388170 457094 388226
rect 457150 388170 457218 388226
rect 457274 388170 457342 388226
rect 457398 388170 457494 388226
rect 456874 388102 457494 388170
rect 456874 388046 456970 388102
rect 457026 388046 457094 388102
rect 457150 388046 457218 388102
rect 457274 388046 457342 388102
rect 457398 388046 457494 388102
rect 456874 387978 457494 388046
rect 456874 387922 456970 387978
rect 457026 387922 457094 387978
rect 457150 387922 457218 387978
rect 457274 387922 457342 387978
rect 457398 387922 457494 387978
rect 456874 370350 457494 387922
rect 456874 370294 456970 370350
rect 457026 370294 457094 370350
rect 457150 370294 457218 370350
rect 457274 370294 457342 370350
rect 457398 370294 457494 370350
rect 456874 370226 457494 370294
rect 456874 370170 456970 370226
rect 457026 370170 457094 370226
rect 457150 370170 457218 370226
rect 457274 370170 457342 370226
rect 457398 370170 457494 370226
rect 456874 370102 457494 370170
rect 456874 370046 456970 370102
rect 457026 370046 457094 370102
rect 457150 370046 457218 370102
rect 457274 370046 457342 370102
rect 457398 370046 457494 370102
rect 456874 369978 457494 370046
rect 456874 369922 456970 369978
rect 457026 369922 457094 369978
rect 457150 369922 457218 369978
rect 457274 369922 457342 369978
rect 457398 369922 457494 369978
rect 456874 352350 457494 369922
rect 456874 352294 456970 352350
rect 457026 352294 457094 352350
rect 457150 352294 457218 352350
rect 457274 352294 457342 352350
rect 457398 352294 457494 352350
rect 456874 352226 457494 352294
rect 456874 352170 456970 352226
rect 457026 352170 457094 352226
rect 457150 352170 457218 352226
rect 457274 352170 457342 352226
rect 457398 352170 457494 352226
rect 456874 352102 457494 352170
rect 456874 352046 456970 352102
rect 457026 352046 457094 352102
rect 457150 352046 457218 352102
rect 457274 352046 457342 352102
rect 457398 352046 457494 352102
rect 456874 351978 457494 352046
rect 456874 351922 456970 351978
rect 457026 351922 457094 351978
rect 457150 351922 457218 351978
rect 457274 351922 457342 351978
rect 457398 351922 457494 351978
rect 456874 334350 457494 351922
rect 456874 334294 456970 334350
rect 457026 334294 457094 334350
rect 457150 334294 457218 334350
rect 457274 334294 457342 334350
rect 457398 334294 457494 334350
rect 456874 334226 457494 334294
rect 456874 334170 456970 334226
rect 457026 334170 457094 334226
rect 457150 334170 457218 334226
rect 457274 334170 457342 334226
rect 457398 334170 457494 334226
rect 456874 334102 457494 334170
rect 456874 334046 456970 334102
rect 457026 334046 457094 334102
rect 457150 334046 457218 334102
rect 457274 334046 457342 334102
rect 457398 334046 457494 334102
rect 456874 333978 457494 334046
rect 456874 333922 456970 333978
rect 457026 333922 457094 333978
rect 457150 333922 457218 333978
rect 457274 333922 457342 333978
rect 457398 333922 457494 333978
rect 456874 316350 457494 333922
rect 456874 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 457494 316350
rect 456874 316226 457494 316294
rect 456874 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 457494 316226
rect 456874 316102 457494 316170
rect 456874 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 457494 316102
rect 456874 315978 457494 316046
rect 456874 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 457494 315978
rect 456874 298350 457494 315922
rect 456874 298294 456970 298350
rect 457026 298294 457094 298350
rect 457150 298294 457218 298350
rect 457274 298294 457342 298350
rect 457398 298294 457494 298350
rect 456874 298226 457494 298294
rect 456874 298170 456970 298226
rect 457026 298170 457094 298226
rect 457150 298170 457218 298226
rect 457274 298170 457342 298226
rect 457398 298170 457494 298226
rect 456874 298102 457494 298170
rect 456874 298046 456970 298102
rect 457026 298046 457094 298102
rect 457150 298046 457218 298102
rect 457274 298046 457342 298102
rect 457398 298046 457494 298102
rect 456874 297978 457494 298046
rect 456874 297922 456970 297978
rect 457026 297922 457094 297978
rect 457150 297922 457218 297978
rect 457274 297922 457342 297978
rect 457398 297922 457494 297978
rect 456874 280350 457494 297922
rect 456874 280294 456970 280350
rect 457026 280294 457094 280350
rect 457150 280294 457218 280350
rect 457274 280294 457342 280350
rect 457398 280294 457494 280350
rect 456874 280226 457494 280294
rect 456874 280170 456970 280226
rect 457026 280170 457094 280226
rect 457150 280170 457218 280226
rect 457274 280170 457342 280226
rect 457398 280170 457494 280226
rect 456874 280102 457494 280170
rect 456874 280046 456970 280102
rect 457026 280046 457094 280102
rect 457150 280046 457218 280102
rect 457274 280046 457342 280102
rect 457398 280046 457494 280102
rect 456874 279978 457494 280046
rect 456874 279922 456970 279978
rect 457026 279922 457094 279978
rect 457150 279922 457218 279978
rect 457274 279922 457342 279978
rect 457398 279922 457494 279978
rect 456874 262350 457494 279922
rect 456874 262294 456970 262350
rect 457026 262294 457094 262350
rect 457150 262294 457218 262350
rect 457274 262294 457342 262350
rect 457398 262294 457494 262350
rect 456874 262226 457494 262294
rect 456874 262170 456970 262226
rect 457026 262170 457094 262226
rect 457150 262170 457218 262226
rect 457274 262170 457342 262226
rect 457398 262170 457494 262226
rect 456874 262102 457494 262170
rect 456874 262046 456970 262102
rect 457026 262046 457094 262102
rect 457150 262046 457218 262102
rect 457274 262046 457342 262102
rect 457398 262046 457494 262102
rect 456874 261978 457494 262046
rect 456874 261922 456970 261978
rect 457026 261922 457094 261978
rect 457150 261922 457218 261978
rect 457274 261922 457342 261978
rect 457398 261922 457494 261978
rect 456874 244350 457494 261922
rect 456874 244294 456970 244350
rect 457026 244294 457094 244350
rect 457150 244294 457218 244350
rect 457274 244294 457342 244350
rect 457398 244294 457494 244350
rect 456874 244226 457494 244294
rect 456874 244170 456970 244226
rect 457026 244170 457094 244226
rect 457150 244170 457218 244226
rect 457274 244170 457342 244226
rect 457398 244170 457494 244226
rect 456874 244102 457494 244170
rect 456874 244046 456970 244102
rect 457026 244046 457094 244102
rect 457150 244046 457218 244102
rect 457274 244046 457342 244102
rect 457398 244046 457494 244102
rect 456874 243978 457494 244046
rect 456874 243922 456970 243978
rect 457026 243922 457094 243978
rect 457150 243922 457218 243978
rect 457274 243922 457342 243978
rect 457398 243922 457494 243978
rect 456874 226350 457494 243922
rect 456874 226294 456970 226350
rect 457026 226294 457094 226350
rect 457150 226294 457218 226350
rect 457274 226294 457342 226350
rect 457398 226294 457494 226350
rect 456874 226226 457494 226294
rect 456874 226170 456970 226226
rect 457026 226170 457094 226226
rect 457150 226170 457218 226226
rect 457274 226170 457342 226226
rect 457398 226170 457494 226226
rect 456874 226102 457494 226170
rect 456874 226046 456970 226102
rect 457026 226046 457094 226102
rect 457150 226046 457218 226102
rect 457274 226046 457342 226102
rect 457398 226046 457494 226102
rect 456874 225978 457494 226046
rect 456874 225922 456970 225978
rect 457026 225922 457094 225978
rect 457150 225922 457218 225978
rect 457274 225922 457342 225978
rect 457398 225922 457494 225978
rect 456874 208350 457494 225922
rect 456874 208294 456970 208350
rect 457026 208294 457094 208350
rect 457150 208294 457218 208350
rect 457274 208294 457342 208350
rect 457398 208294 457494 208350
rect 456874 208226 457494 208294
rect 456874 208170 456970 208226
rect 457026 208170 457094 208226
rect 457150 208170 457218 208226
rect 457274 208170 457342 208226
rect 457398 208170 457494 208226
rect 456874 208102 457494 208170
rect 456874 208046 456970 208102
rect 457026 208046 457094 208102
rect 457150 208046 457218 208102
rect 457274 208046 457342 208102
rect 457398 208046 457494 208102
rect 456874 207978 457494 208046
rect 456874 207922 456970 207978
rect 457026 207922 457094 207978
rect 457150 207922 457218 207978
rect 457274 207922 457342 207978
rect 457398 207922 457494 207978
rect 456874 190350 457494 207922
rect 456874 190294 456970 190350
rect 457026 190294 457094 190350
rect 457150 190294 457218 190350
rect 457274 190294 457342 190350
rect 457398 190294 457494 190350
rect 456874 190226 457494 190294
rect 456874 190170 456970 190226
rect 457026 190170 457094 190226
rect 457150 190170 457218 190226
rect 457274 190170 457342 190226
rect 457398 190170 457494 190226
rect 456874 190102 457494 190170
rect 456874 190046 456970 190102
rect 457026 190046 457094 190102
rect 457150 190046 457218 190102
rect 457274 190046 457342 190102
rect 457398 190046 457494 190102
rect 456874 189978 457494 190046
rect 456874 189922 456970 189978
rect 457026 189922 457094 189978
rect 457150 189922 457218 189978
rect 457274 189922 457342 189978
rect 457398 189922 457494 189978
rect 456874 172350 457494 189922
rect 456874 172294 456970 172350
rect 457026 172294 457094 172350
rect 457150 172294 457218 172350
rect 457274 172294 457342 172350
rect 457398 172294 457494 172350
rect 456874 172226 457494 172294
rect 456874 172170 456970 172226
rect 457026 172170 457094 172226
rect 457150 172170 457218 172226
rect 457274 172170 457342 172226
rect 457398 172170 457494 172226
rect 456874 172102 457494 172170
rect 456874 172046 456970 172102
rect 457026 172046 457094 172102
rect 457150 172046 457218 172102
rect 457274 172046 457342 172102
rect 457398 172046 457494 172102
rect 456874 171978 457494 172046
rect 456874 171922 456970 171978
rect 457026 171922 457094 171978
rect 457150 171922 457218 171978
rect 457274 171922 457342 171978
rect 457398 171922 457494 171978
rect 456874 154350 457494 171922
rect 456874 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 457494 154350
rect 456874 154226 457494 154294
rect 456874 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 457494 154226
rect 456874 154102 457494 154170
rect 456874 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 457494 154102
rect 456874 153978 457494 154046
rect 456874 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 457494 153978
rect 456874 136350 457494 153922
rect 456874 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 457494 136350
rect 456874 136226 457494 136294
rect 456874 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 457494 136226
rect 456874 136102 457494 136170
rect 456874 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 457494 136102
rect 456874 135978 457494 136046
rect 456874 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 457494 135978
rect 456874 118350 457494 135922
rect 456874 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 457494 118350
rect 456874 118226 457494 118294
rect 456874 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 457494 118226
rect 456874 118102 457494 118170
rect 456874 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 457494 118102
rect 456874 117978 457494 118046
rect 456874 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 457494 117978
rect 456874 100350 457494 117922
rect 456874 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 457494 100350
rect 456874 100226 457494 100294
rect 456874 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 457494 100226
rect 456874 100102 457494 100170
rect 456874 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 457494 100102
rect 456874 99978 457494 100046
rect 456874 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 457494 99978
rect 456874 82350 457494 99922
rect 456874 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 457494 82350
rect 456874 82226 457494 82294
rect 456874 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 457494 82226
rect 456874 82102 457494 82170
rect 456874 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 457494 82102
rect 456874 81978 457494 82046
rect 456874 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 457494 81978
rect 456874 64350 457494 81922
rect 456874 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 457494 64350
rect 456874 64226 457494 64294
rect 456874 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 457494 64226
rect 456874 64102 457494 64170
rect 456874 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 457494 64102
rect 456874 63978 457494 64046
rect 456874 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 457494 63978
rect 456874 46350 457494 63922
rect 456874 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 457494 46350
rect 456874 46226 457494 46294
rect 456874 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 457494 46226
rect 456874 46102 457494 46170
rect 456874 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 457494 46102
rect 456874 45978 457494 46046
rect 456874 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 457494 45978
rect 456874 28350 457494 45922
rect 456874 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 457494 28350
rect 456874 28226 457494 28294
rect 456874 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 457494 28226
rect 456874 28102 457494 28170
rect 456874 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 457494 28102
rect 456874 27978 457494 28046
rect 456874 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 457494 27978
rect 456874 10350 457494 27922
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 526350 471774 543922
rect 471154 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 471774 526350
rect 471154 526226 471774 526294
rect 471154 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 471774 526226
rect 471154 526102 471774 526170
rect 471154 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 471774 526102
rect 471154 525978 471774 526046
rect 471154 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 471774 525978
rect 471154 508350 471774 525922
rect 471154 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 471774 508350
rect 471154 508226 471774 508294
rect 471154 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 471774 508226
rect 471154 508102 471774 508170
rect 471154 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 471774 508102
rect 471154 507978 471774 508046
rect 471154 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 471774 507978
rect 471154 490350 471774 507922
rect 471154 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 471774 490350
rect 471154 490226 471774 490294
rect 471154 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 471774 490226
rect 471154 490102 471774 490170
rect 471154 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 471774 490102
rect 471154 489978 471774 490046
rect 471154 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 471774 489978
rect 471154 472350 471774 489922
rect 471154 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 471774 472350
rect 471154 472226 471774 472294
rect 471154 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 471774 472226
rect 471154 472102 471774 472170
rect 471154 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 471774 472102
rect 471154 471978 471774 472046
rect 471154 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 471774 471978
rect 471154 454350 471774 471922
rect 471154 454294 471250 454350
rect 471306 454294 471374 454350
rect 471430 454294 471498 454350
rect 471554 454294 471622 454350
rect 471678 454294 471774 454350
rect 471154 454226 471774 454294
rect 471154 454170 471250 454226
rect 471306 454170 471374 454226
rect 471430 454170 471498 454226
rect 471554 454170 471622 454226
rect 471678 454170 471774 454226
rect 471154 454102 471774 454170
rect 471154 454046 471250 454102
rect 471306 454046 471374 454102
rect 471430 454046 471498 454102
rect 471554 454046 471622 454102
rect 471678 454046 471774 454102
rect 471154 453978 471774 454046
rect 471154 453922 471250 453978
rect 471306 453922 471374 453978
rect 471430 453922 471498 453978
rect 471554 453922 471622 453978
rect 471678 453922 471774 453978
rect 471154 436350 471774 453922
rect 471154 436294 471250 436350
rect 471306 436294 471374 436350
rect 471430 436294 471498 436350
rect 471554 436294 471622 436350
rect 471678 436294 471774 436350
rect 471154 436226 471774 436294
rect 471154 436170 471250 436226
rect 471306 436170 471374 436226
rect 471430 436170 471498 436226
rect 471554 436170 471622 436226
rect 471678 436170 471774 436226
rect 471154 436102 471774 436170
rect 471154 436046 471250 436102
rect 471306 436046 471374 436102
rect 471430 436046 471498 436102
rect 471554 436046 471622 436102
rect 471678 436046 471774 436102
rect 471154 435978 471774 436046
rect 471154 435922 471250 435978
rect 471306 435922 471374 435978
rect 471430 435922 471498 435978
rect 471554 435922 471622 435978
rect 471678 435922 471774 435978
rect 471154 418350 471774 435922
rect 471154 418294 471250 418350
rect 471306 418294 471374 418350
rect 471430 418294 471498 418350
rect 471554 418294 471622 418350
rect 471678 418294 471774 418350
rect 471154 418226 471774 418294
rect 471154 418170 471250 418226
rect 471306 418170 471374 418226
rect 471430 418170 471498 418226
rect 471554 418170 471622 418226
rect 471678 418170 471774 418226
rect 471154 418102 471774 418170
rect 471154 418046 471250 418102
rect 471306 418046 471374 418102
rect 471430 418046 471498 418102
rect 471554 418046 471622 418102
rect 471678 418046 471774 418102
rect 471154 417978 471774 418046
rect 471154 417922 471250 417978
rect 471306 417922 471374 417978
rect 471430 417922 471498 417978
rect 471554 417922 471622 417978
rect 471678 417922 471774 417978
rect 471154 400350 471774 417922
rect 471154 400294 471250 400350
rect 471306 400294 471374 400350
rect 471430 400294 471498 400350
rect 471554 400294 471622 400350
rect 471678 400294 471774 400350
rect 471154 400226 471774 400294
rect 471154 400170 471250 400226
rect 471306 400170 471374 400226
rect 471430 400170 471498 400226
rect 471554 400170 471622 400226
rect 471678 400170 471774 400226
rect 471154 400102 471774 400170
rect 471154 400046 471250 400102
rect 471306 400046 471374 400102
rect 471430 400046 471498 400102
rect 471554 400046 471622 400102
rect 471678 400046 471774 400102
rect 471154 399978 471774 400046
rect 471154 399922 471250 399978
rect 471306 399922 471374 399978
rect 471430 399922 471498 399978
rect 471554 399922 471622 399978
rect 471678 399922 471774 399978
rect 471154 382350 471774 399922
rect 471154 382294 471250 382350
rect 471306 382294 471374 382350
rect 471430 382294 471498 382350
rect 471554 382294 471622 382350
rect 471678 382294 471774 382350
rect 471154 382226 471774 382294
rect 471154 382170 471250 382226
rect 471306 382170 471374 382226
rect 471430 382170 471498 382226
rect 471554 382170 471622 382226
rect 471678 382170 471774 382226
rect 471154 382102 471774 382170
rect 471154 382046 471250 382102
rect 471306 382046 471374 382102
rect 471430 382046 471498 382102
rect 471554 382046 471622 382102
rect 471678 382046 471774 382102
rect 471154 381978 471774 382046
rect 471154 381922 471250 381978
rect 471306 381922 471374 381978
rect 471430 381922 471498 381978
rect 471554 381922 471622 381978
rect 471678 381922 471774 381978
rect 471154 364350 471774 381922
rect 471154 364294 471250 364350
rect 471306 364294 471374 364350
rect 471430 364294 471498 364350
rect 471554 364294 471622 364350
rect 471678 364294 471774 364350
rect 471154 364226 471774 364294
rect 471154 364170 471250 364226
rect 471306 364170 471374 364226
rect 471430 364170 471498 364226
rect 471554 364170 471622 364226
rect 471678 364170 471774 364226
rect 471154 364102 471774 364170
rect 471154 364046 471250 364102
rect 471306 364046 471374 364102
rect 471430 364046 471498 364102
rect 471554 364046 471622 364102
rect 471678 364046 471774 364102
rect 471154 363978 471774 364046
rect 471154 363922 471250 363978
rect 471306 363922 471374 363978
rect 471430 363922 471498 363978
rect 471554 363922 471622 363978
rect 471678 363922 471774 363978
rect 471154 346350 471774 363922
rect 471154 346294 471250 346350
rect 471306 346294 471374 346350
rect 471430 346294 471498 346350
rect 471554 346294 471622 346350
rect 471678 346294 471774 346350
rect 471154 346226 471774 346294
rect 471154 346170 471250 346226
rect 471306 346170 471374 346226
rect 471430 346170 471498 346226
rect 471554 346170 471622 346226
rect 471678 346170 471774 346226
rect 471154 346102 471774 346170
rect 471154 346046 471250 346102
rect 471306 346046 471374 346102
rect 471430 346046 471498 346102
rect 471554 346046 471622 346102
rect 471678 346046 471774 346102
rect 471154 345978 471774 346046
rect 471154 345922 471250 345978
rect 471306 345922 471374 345978
rect 471430 345922 471498 345978
rect 471554 345922 471622 345978
rect 471678 345922 471774 345978
rect 471154 328350 471774 345922
rect 471154 328294 471250 328350
rect 471306 328294 471374 328350
rect 471430 328294 471498 328350
rect 471554 328294 471622 328350
rect 471678 328294 471774 328350
rect 471154 328226 471774 328294
rect 471154 328170 471250 328226
rect 471306 328170 471374 328226
rect 471430 328170 471498 328226
rect 471554 328170 471622 328226
rect 471678 328170 471774 328226
rect 471154 328102 471774 328170
rect 471154 328046 471250 328102
rect 471306 328046 471374 328102
rect 471430 328046 471498 328102
rect 471554 328046 471622 328102
rect 471678 328046 471774 328102
rect 471154 327978 471774 328046
rect 471154 327922 471250 327978
rect 471306 327922 471374 327978
rect 471430 327922 471498 327978
rect 471554 327922 471622 327978
rect 471678 327922 471774 327978
rect 471154 310350 471774 327922
rect 471154 310294 471250 310350
rect 471306 310294 471374 310350
rect 471430 310294 471498 310350
rect 471554 310294 471622 310350
rect 471678 310294 471774 310350
rect 471154 310226 471774 310294
rect 471154 310170 471250 310226
rect 471306 310170 471374 310226
rect 471430 310170 471498 310226
rect 471554 310170 471622 310226
rect 471678 310170 471774 310226
rect 471154 310102 471774 310170
rect 471154 310046 471250 310102
rect 471306 310046 471374 310102
rect 471430 310046 471498 310102
rect 471554 310046 471622 310102
rect 471678 310046 471774 310102
rect 471154 309978 471774 310046
rect 471154 309922 471250 309978
rect 471306 309922 471374 309978
rect 471430 309922 471498 309978
rect 471554 309922 471622 309978
rect 471678 309922 471774 309978
rect 471154 292350 471774 309922
rect 471154 292294 471250 292350
rect 471306 292294 471374 292350
rect 471430 292294 471498 292350
rect 471554 292294 471622 292350
rect 471678 292294 471774 292350
rect 471154 292226 471774 292294
rect 471154 292170 471250 292226
rect 471306 292170 471374 292226
rect 471430 292170 471498 292226
rect 471554 292170 471622 292226
rect 471678 292170 471774 292226
rect 471154 292102 471774 292170
rect 471154 292046 471250 292102
rect 471306 292046 471374 292102
rect 471430 292046 471498 292102
rect 471554 292046 471622 292102
rect 471678 292046 471774 292102
rect 471154 291978 471774 292046
rect 471154 291922 471250 291978
rect 471306 291922 471374 291978
rect 471430 291922 471498 291978
rect 471554 291922 471622 291978
rect 471678 291922 471774 291978
rect 471154 274350 471774 291922
rect 471154 274294 471250 274350
rect 471306 274294 471374 274350
rect 471430 274294 471498 274350
rect 471554 274294 471622 274350
rect 471678 274294 471774 274350
rect 471154 274226 471774 274294
rect 471154 274170 471250 274226
rect 471306 274170 471374 274226
rect 471430 274170 471498 274226
rect 471554 274170 471622 274226
rect 471678 274170 471774 274226
rect 471154 274102 471774 274170
rect 471154 274046 471250 274102
rect 471306 274046 471374 274102
rect 471430 274046 471498 274102
rect 471554 274046 471622 274102
rect 471678 274046 471774 274102
rect 471154 273978 471774 274046
rect 471154 273922 471250 273978
rect 471306 273922 471374 273978
rect 471430 273922 471498 273978
rect 471554 273922 471622 273978
rect 471678 273922 471774 273978
rect 471154 256350 471774 273922
rect 471154 256294 471250 256350
rect 471306 256294 471374 256350
rect 471430 256294 471498 256350
rect 471554 256294 471622 256350
rect 471678 256294 471774 256350
rect 471154 256226 471774 256294
rect 471154 256170 471250 256226
rect 471306 256170 471374 256226
rect 471430 256170 471498 256226
rect 471554 256170 471622 256226
rect 471678 256170 471774 256226
rect 471154 256102 471774 256170
rect 471154 256046 471250 256102
rect 471306 256046 471374 256102
rect 471430 256046 471498 256102
rect 471554 256046 471622 256102
rect 471678 256046 471774 256102
rect 471154 255978 471774 256046
rect 471154 255922 471250 255978
rect 471306 255922 471374 255978
rect 471430 255922 471498 255978
rect 471554 255922 471622 255978
rect 471678 255922 471774 255978
rect 471154 238350 471774 255922
rect 471154 238294 471250 238350
rect 471306 238294 471374 238350
rect 471430 238294 471498 238350
rect 471554 238294 471622 238350
rect 471678 238294 471774 238350
rect 471154 238226 471774 238294
rect 471154 238170 471250 238226
rect 471306 238170 471374 238226
rect 471430 238170 471498 238226
rect 471554 238170 471622 238226
rect 471678 238170 471774 238226
rect 471154 238102 471774 238170
rect 471154 238046 471250 238102
rect 471306 238046 471374 238102
rect 471430 238046 471498 238102
rect 471554 238046 471622 238102
rect 471678 238046 471774 238102
rect 471154 237978 471774 238046
rect 471154 237922 471250 237978
rect 471306 237922 471374 237978
rect 471430 237922 471498 237978
rect 471554 237922 471622 237978
rect 471678 237922 471774 237978
rect 471154 220350 471774 237922
rect 471154 220294 471250 220350
rect 471306 220294 471374 220350
rect 471430 220294 471498 220350
rect 471554 220294 471622 220350
rect 471678 220294 471774 220350
rect 471154 220226 471774 220294
rect 471154 220170 471250 220226
rect 471306 220170 471374 220226
rect 471430 220170 471498 220226
rect 471554 220170 471622 220226
rect 471678 220170 471774 220226
rect 471154 220102 471774 220170
rect 471154 220046 471250 220102
rect 471306 220046 471374 220102
rect 471430 220046 471498 220102
rect 471554 220046 471622 220102
rect 471678 220046 471774 220102
rect 471154 219978 471774 220046
rect 471154 219922 471250 219978
rect 471306 219922 471374 219978
rect 471430 219922 471498 219978
rect 471554 219922 471622 219978
rect 471678 219922 471774 219978
rect 471154 202350 471774 219922
rect 471154 202294 471250 202350
rect 471306 202294 471374 202350
rect 471430 202294 471498 202350
rect 471554 202294 471622 202350
rect 471678 202294 471774 202350
rect 471154 202226 471774 202294
rect 471154 202170 471250 202226
rect 471306 202170 471374 202226
rect 471430 202170 471498 202226
rect 471554 202170 471622 202226
rect 471678 202170 471774 202226
rect 471154 202102 471774 202170
rect 471154 202046 471250 202102
rect 471306 202046 471374 202102
rect 471430 202046 471498 202102
rect 471554 202046 471622 202102
rect 471678 202046 471774 202102
rect 471154 201978 471774 202046
rect 471154 201922 471250 201978
rect 471306 201922 471374 201978
rect 471430 201922 471498 201978
rect 471554 201922 471622 201978
rect 471678 201922 471774 201978
rect 471154 184350 471774 201922
rect 471154 184294 471250 184350
rect 471306 184294 471374 184350
rect 471430 184294 471498 184350
rect 471554 184294 471622 184350
rect 471678 184294 471774 184350
rect 471154 184226 471774 184294
rect 471154 184170 471250 184226
rect 471306 184170 471374 184226
rect 471430 184170 471498 184226
rect 471554 184170 471622 184226
rect 471678 184170 471774 184226
rect 471154 184102 471774 184170
rect 471154 184046 471250 184102
rect 471306 184046 471374 184102
rect 471430 184046 471498 184102
rect 471554 184046 471622 184102
rect 471678 184046 471774 184102
rect 471154 183978 471774 184046
rect 471154 183922 471250 183978
rect 471306 183922 471374 183978
rect 471430 183922 471498 183978
rect 471554 183922 471622 183978
rect 471678 183922 471774 183978
rect 471154 166350 471774 183922
rect 471154 166294 471250 166350
rect 471306 166294 471374 166350
rect 471430 166294 471498 166350
rect 471554 166294 471622 166350
rect 471678 166294 471774 166350
rect 471154 166226 471774 166294
rect 471154 166170 471250 166226
rect 471306 166170 471374 166226
rect 471430 166170 471498 166226
rect 471554 166170 471622 166226
rect 471678 166170 471774 166226
rect 471154 166102 471774 166170
rect 471154 166046 471250 166102
rect 471306 166046 471374 166102
rect 471430 166046 471498 166102
rect 471554 166046 471622 166102
rect 471678 166046 471774 166102
rect 471154 165978 471774 166046
rect 471154 165922 471250 165978
rect 471306 165922 471374 165978
rect 471430 165922 471498 165978
rect 471554 165922 471622 165978
rect 471678 165922 471774 165978
rect 471154 148350 471774 165922
rect 471154 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 471774 148350
rect 471154 148226 471774 148294
rect 471154 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 471774 148226
rect 471154 148102 471774 148170
rect 471154 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 471774 148102
rect 471154 147978 471774 148046
rect 471154 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 471774 147978
rect 471154 130350 471774 147922
rect 471154 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 471774 130350
rect 471154 130226 471774 130294
rect 471154 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 471774 130226
rect 471154 130102 471774 130170
rect 471154 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 471774 130102
rect 471154 129978 471774 130046
rect 471154 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 471774 129978
rect 471154 112350 471774 129922
rect 471154 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 471774 112350
rect 471154 112226 471774 112294
rect 471154 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 471774 112226
rect 471154 112102 471774 112170
rect 471154 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 471774 112102
rect 471154 111978 471774 112046
rect 471154 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 471774 111978
rect 471154 94350 471774 111922
rect 471154 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 471774 94350
rect 471154 94226 471774 94294
rect 471154 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 471774 94226
rect 471154 94102 471774 94170
rect 471154 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 471774 94102
rect 471154 93978 471774 94046
rect 471154 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 471774 93978
rect 471154 76350 471774 93922
rect 471154 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 471774 76350
rect 471154 76226 471774 76294
rect 471154 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 471774 76226
rect 471154 76102 471774 76170
rect 471154 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 471774 76102
rect 471154 75978 471774 76046
rect 471154 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 471774 75978
rect 471154 58350 471774 75922
rect 471154 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 471774 58350
rect 471154 58226 471774 58294
rect 471154 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 471774 58226
rect 471154 58102 471774 58170
rect 471154 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 471774 58102
rect 471154 57978 471774 58046
rect 471154 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 471774 57978
rect 471154 40350 471774 57922
rect 471154 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 471774 40350
rect 471154 40226 471774 40294
rect 471154 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 471774 40226
rect 471154 40102 471774 40170
rect 471154 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 471774 40102
rect 471154 39978 471774 40046
rect 471154 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 471774 39978
rect 471154 22350 471774 39922
rect 471154 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 471774 22350
rect 471154 22226 471774 22294
rect 471154 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 471774 22226
rect 471154 22102 471774 22170
rect 471154 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 471774 22102
rect 471154 21978 471774 22046
rect 471154 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 471774 21978
rect 471154 4350 471774 21922
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 598172 475494 598268
rect 474874 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 475494 598172
rect 474874 598048 475494 598116
rect 474874 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 475494 598048
rect 474874 597924 475494 597992
rect 474874 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 475494 597924
rect 474874 597800 475494 597868
rect 474874 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 475494 597800
rect 474874 586350 475494 597744
rect 474874 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 475494 586350
rect 474874 586226 475494 586294
rect 474874 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 475494 586226
rect 474874 586102 475494 586170
rect 474874 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 475494 586102
rect 474874 585978 475494 586046
rect 474874 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 475494 585978
rect 474874 568350 475494 585922
rect 474874 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 475494 568350
rect 474874 568226 475494 568294
rect 474874 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 475494 568226
rect 474874 568102 475494 568170
rect 474874 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 475494 568102
rect 474874 567978 475494 568046
rect 474874 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 475494 567978
rect 474874 550350 475494 567922
rect 474874 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 475494 550350
rect 474874 550226 475494 550294
rect 474874 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 475494 550226
rect 474874 550102 475494 550170
rect 474874 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 475494 550102
rect 474874 549978 475494 550046
rect 474874 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 475494 549978
rect 474874 532350 475494 549922
rect 474874 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 475494 532350
rect 474874 532226 475494 532294
rect 474874 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 475494 532226
rect 474874 532102 475494 532170
rect 474874 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 475494 532102
rect 474874 531978 475494 532046
rect 474874 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 475494 531978
rect 474874 514350 475494 531922
rect 474874 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 475494 514350
rect 474874 514226 475494 514294
rect 474874 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 475494 514226
rect 474874 514102 475494 514170
rect 474874 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 475494 514102
rect 474874 513978 475494 514046
rect 474874 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 475494 513978
rect 474874 496350 475494 513922
rect 474874 496294 474970 496350
rect 475026 496294 475094 496350
rect 475150 496294 475218 496350
rect 475274 496294 475342 496350
rect 475398 496294 475494 496350
rect 474874 496226 475494 496294
rect 474874 496170 474970 496226
rect 475026 496170 475094 496226
rect 475150 496170 475218 496226
rect 475274 496170 475342 496226
rect 475398 496170 475494 496226
rect 474874 496102 475494 496170
rect 474874 496046 474970 496102
rect 475026 496046 475094 496102
rect 475150 496046 475218 496102
rect 475274 496046 475342 496102
rect 475398 496046 475494 496102
rect 474874 495978 475494 496046
rect 474874 495922 474970 495978
rect 475026 495922 475094 495978
rect 475150 495922 475218 495978
rect 475274 495922 475342 495978
rect 475398 495922 475494 495978
rect 474874 478350 475494 495922
rect 474874 478294 474970 478350
rect 475026 478294 475094 478350
rect 475150 478294 475218 478350
rect 475274 478294 475342 478350
rect 475398 478294 475494 478350
rect 474874 478226 475494 478294
rect 474874 478170 474970 478226
rect 475026 478170 475094 478226
rect 475150 478170 475218 478226
rect 475274 478170 475342 478226
rect 475398 478170 475494 478226
rect 474874 478102 475494 478170
rect 474874 478046 474970 478102
rect 475026 478046 475094 478102
rect 475150 478046 475218 478102
rect 475274 478046 475342 478102
rect 475398 478046 475494 478102
rect 474874 477978 475494 478046
rect 474874 477922 474970 477978
rect 475026 477922 475094 477978
rect 475150 477922 475218 477978
rect 475274 477922 475342 477978
rect 475398 477922 475494 477978
rect 474874 460350 475494 477922
rect 474874 460294 474970 460350
rect 475026 460294 475094 460350
rect 475150 460294 475218 460350
rect 475274 460294 475342 460350
rect 475398 460294 475494 460350
rect 474874 460226 475494 460294
rect 474874 460170 474970 460226
rect 475026 460170 475094 460226
rect 475150 460170 475218 460226
rect 475274 460170 475342 460226
rect 475398 460170 475494 460226
rect 474874 460102 475494 460170
rect 474874 460046 474970 460102
rect 475026 460046 475094 460102
rect 475150 460046 475218 460102
rect 475274 460046 475342 460102
rect 475398 460046 475494 460102
rect 474874 459978 475494 460046
rect 474874 459922 474970 459978
rect 475026 459922 475094 459978
rect 475150 459922 475218 459978
rect 475274 459922 475342 459978
rect 475398 459922 475494 459978
rect 474874 442350 475494 459922
rect 474874 442294 474970 442350
rect 475026 442294 475094 442350
rect 475150 442294 475218 442350
rect 475274 442294 475342 442350
rect 475398 442294 475494 442350
rect 474874 442226 475494 442294
rect 474874 442170 474970 442226
rect 475026 442170 475094 442226
rect 475150 442170 475218 442226
rect 475274 442170 475342 442226
rect 475398 442170 475494 442226
rect 474874 442102 475494 442170
rect 474874 442046 474970 442102
rect 475026 442046 475094 442102
rect 475150 442046 475218 442102
rect 475274 442046 475342 442102
rect 475398 442046 475494 442102
rect 474874 441978 475494 442046
rect 474874 441922 474970 441978
rect 475026 441922 475094 441978
rect 475150 441922 475218 441978
rect 475274 441922 475342 441978
rect 475398 441922 475494 441978
rect 474874 424350 475494 441922
rect 474874 424294 474970 424350
rect 475026 424294 475094 424350
rect 475150 424294 475218 424350
rect 475274 424294 475342 424350
rect 475398 424294 475494 424350
rect 474874 424226 475494 424294
rect 474874 424170 474970 424226
rect 475026 424170 475094 424226
rect 475150 424170 475218 424226
rect 475274 424170 475342 424226
rect 475398 424170 475494 424226
rect 474874 424102 475494 424170
rect 474874 424046 474970 424102
rect 475026 424046 475094 424102
rect 475150 424046 475218 424102
rect 475274 424046 475342 424102
rect 475398 424046 475494 424102
rect 474874 423978 475494 424046
rect 474874 423922 474970 423978
rect 475026 423922 475094 423978
rect 475150 423922 475218 423978
rect 475274 423922 475342 423978
rect 475398 423922 475494 423978
rect 474874 406350 475494 423922
rect 474874 406294 474970 406350
rect 475026 406294 475094 406350
rect 475150 406294 475218 406350
rect 475274 406294 475342 406350
rect 475398 406294 475494 406350
rect 474874 406226 475494 406294
rect 474874 406170 474970 406226
rect 475026 406170 475094 406226
rect 475150 406170 475218 406226
rect 475274 406170 475342 406226
rect 475398 406170 475494 406226
rect 474874 406102 475494 406170
rect 474874 406046 474970 406102
rect 475026 406046 475094 406102
rect 475150 406046 475218 406102
rect 475274 406046 475342 406102
rect 475398 406046 475494 406102
rect 474874 405978 475494 406046
rect 474874 405922 474970 405978
rect 475026 405922 475094 405978
rect 475150 405922 475218 405978
rect 475274 405922 475342 405978
rect 475398 405922 475494 405978
rect 474874 388350 475494 405922
rect 474874 388294 474970 388350
rect 475026 388294 475094 388350
rect 475150 388294 475218 388350
rect 475274 388294 475342 388350
rect 475398 388294 475494 388350
rect 474874 388226 475494 388294
rect 474874 388170 474970 388226
rect 475026 388170 475094 388226
rect 475150 388170 475218 388226
rect 475274 388170 475342 388226
rect 475398 388170 475494 388226
rect 474874 388102 475494 388170
rect 474874 388046 474970 388102
rect 475026 388046 475094 388102
rect 475150 388046 475218 388102
rect 475274 388046 475342 388102
rect 475398 388046 475494 388102
rect 474874 387978 475494 388046
rect 474874 387922 474970 387978
rect 475026 387922 475094 387978
rect 475150 387922 475218 387978
rect 475274 387922 475342 387978
rect 475398 387922 475494 387978
rect 474874 370350 475494 387922
rect 474874 370294 474970 370350
rect 475026 370294 475094 370350
rect 475150 370294 475218 370350
rect 475274 370294 475342 370350
rect 475398 370294 475494 370350
rect 474874 370226 475494 370294
rect 474874 370170 474970 370226
rect 475026 370170 475094 370226
rect 475150 370170 475218 370226
rect 475274 370170 475342 370226
rect 475398 370170 475494 370226
rect 474874 370102 475494 370170
rect 474874 370046 474970 370102
rect 475026 370046 475094 370102
rect 475150 370046 475218 370102
rect 475274 370046 475342 370102
rect 475398 370046 475494 370102
rect 474874 369978 475494 370046
rect 474874 369922 474970 369978
rect 475026 369922 475094 369978
rect 475150 369922 475218 369978
rect 475274 369922 475342 369978
rect 475398 369922 475494 369978
rect 474874 352350 475494 369922
rect 474874 352294 474970 352350
rect 475026 352294 475094 352350
rect 475150 352294 475218 352350
rect 475274 352294 475342 352350
rect 475398 352294 475494 352350
rect 474874 352226 475494 352294
rect 474874 352170 474970 352226
rect 475026 352170 475094 352226
rect 475150 352170 475218 352226
rect 475274 352170 475342 352226
rect 475398 352170 475494 352226
rect 474874 352102 475494 352170
rect 474874 352046 474970 352102
rect 475026 352046 475094 352102
rect 475150 352046 475218 352102
rect 475274 352046 475342 352102
rect 475398 352046 475494 352102
rect 474874 351978 475494 352046
rect 474874 351922 474970 351978
rect 475026 351922 475094 351978
rect 475150 351922 475218 351978
rect 475274 351922 475342 351978
rect 475398 351922 475494 351978
rect 474874 334350 475494 351922
rect 474874 334294 474970 334350
rect 475026 334294 475094 334350
rect 475150 334294 475218 334350
rect 475274 334294 475342 334350
rect 475398 334294 475494 334350
rect 474874 334226 475494 334294
rect 474874 334170 474970 334226
rect 475026 334170 475094 334226
rect 475150 334170 475218 334226
rect 475274 334170 475342 334226
rect 475398 334170 475494 334226
rect 474874 334102 475494 334170
rect 474874 334046 474970 334102
rect 475026 334046 475094 334102
rect 475150 334046 475218 334102
rect 475274 334046 475342 334102
rect 475398 334046 475494 334102
rect 474874 333978 475494 334046
rect 474874 333922 474970 333978
rect 475026 333922 475094 333978
rect 475150 333922 475218 333978
rect 475274 333922 475342 333978
rect 475398 333922 475494 333978
rect 474874 316350 475494 333922
rect 474874 316294 474970 316350
rect 475026 316294 475094 316350
rect 475150 316294 475218 316350
rect 475274 316294 475342 316350
rect 475398 316294 475494 316350
rect 474874 316226 475494 316294
rect 474874 316170 474970 316226
rect 475026 316170 475094 316226
rect 475150 316170 475218 316226
rect 475274 316170 475342 316226
rect 475398 316170 475494 316226
rect 474874 316102 475494 316170
rect 474874 316046 474970 316102
rect 475026 316046 475094 316102
rect 475150 316046 475218 316102
rect 475274 316046 475342 316102
rect 475398 316046 475494 316102
rect 474874 315978 475494 316046
rect 474874 315922 474970 315978
rect 475026 315922 475094 315978
rect 475150 315922 475218 315978
rect 475274 315922 475342 315978
rect 475398 315922 475494 315978
rect 474874 298350 475494 315922
rect 474874 298294 474970 298350
rect 475026 298294 475094 298350
rect 475150 298294 475218 298350
rect 475274 298294 475342 298350
rect 475398 298294 475494 298350
rect 474874 298226 475494 298294
rect 474874 298170 474970 298226
rect 475026 298170 475094 298226
rect 475150 298170 475218 298226
rect 475274 298170 475342 298226
rect 475398 298170 475494 298226
rect 474874 298102 475494 298170
rect 474874 298046 474970 298102
rect 475026 298046 475094 298102
rect 475150 298046 475218 298102
rect 475274 298046 475342 298102
rect 475398 298046 475494 298102
rect 474874 297978 475494 298046
rect 474874 297922 474970 297978
rect 475026 297922 475094 297978
rect 475150 297922 475218 297978
rect 475274 297922 475342 297978
rect 475398 297922 475494 297978
rect 474874 280350 475494 297922
rect 474874 280294 474970 280350
rect 475026 280294 475094 280350
rect 475150 280294 475218 280350
rect 475274 280294 475342 280350
rect 475398 280294 475494 280350
rect 474874 280226 475494 280294
rect 474874 280170 474970 280226
rect 475026 280170 475094 280226
rect 475150 280170 475218 280226
rect 475274 280170 475342 280226
rect 475398 280170 475494 280226
rect 474874 280102 475494 280170
rect 474874 280046 474970 280102
rect 475026 280046 475094 280102
rect 475150 280046 475218 280102
rect 475274 280046 475342 280102
rect 475398 280046 475494 280102
rect 474874 279978 475494 280046
rect 474874 279922 474970 279978
rect 475026 279922 475094 279978
rect 475150 279922 475218 279978
rect 475274 279922 475342 279978
rect 475398 279922 475494 279978
rect 474874 262350 475494 279922
rect 474874 262294 474970 262350
rect 475026 262294 475094 262350
rect 475150 262294 475218 262350
rect 475274 262294 475342 262350
rect 475398 262294 475494 262350
rect 474874 262226 475494 262294
rect 474874 262170 474970 262226
rect 475026 262170 475094 262226
rect 475150 262170 475218 262226
rect 475274 262170 475342 262226
rect 475398 262170 475494 262226
rect 474874 262102 475494 262170
rect 474874 262046 474970 262102
rect 475026 262046 475094 262102
rect 475150 262046 475218 262102
rect 475274 262046 475342 262102
rect 475398 262046 475494 262102
rect 474874 261978 475494 262046
rect 474874 261922 474970 261978
rect 475026 261922 475094 261978
rect 475150 261922 475218 261978
rect 475274 261922 475342 261978
rect 475398 261922 475494 261978
rect 474874 244350 475494 261922
rect 474874 244294 474970 244350
rect 475026 244294 475094 244350
rect 475150 244294 475218 244350
rect 475274 244294 475342 244350
rect 475398 244294 475494 244350
rect 474874 244226 475494 244294
rect 474874 244170 474970 244226
rect 475026 244170 475094 244226
rect 475150 244170 475218 244226
rect 475274 244170 475342 244226
rect 475398 244170 475494 244226
rect 474874 244102 475494 244170
rect 474874 244046 474970 244102
rect 475026 244046 475094 244102
rect 475150 244046 475218 244102
rect 475274 244046 475342 244102
rect 475398 244046 475494 244102
rect 474874 243978 475494 244046
rect 474874 243922 474970 243978
rect 475026 243922 475094 243978
rect 475150 243922 475218 243978
rect 475274 243922 475342 243978
rect 475398 243922 475494 243978
rect 474874 226350 475494 243922
rect 474874 226294 474970 226350
rect 475026 226294 475094 226350
rect 475150 226294 475218 226350
rect 475274 226294 475342 226350
rect 475398 226294 475494 226350
rect 474874 226226 475494 226294
rect 474874 226170 474970 226226
rect 475026 226170 475094 226226
rect 475150 226170 475218 226226
rect 475274 226170 475342 226226
rect 475398 226170 475494 226226
rect 474874 226102 475494 226170
rect 474874 226046 474970 226102
rect 475026 226046 475094 226102
rect 475150 226046 475218 226102
rect 475274 226046 475342 226102
rect 475398 226046 475494 226102
rect 474874 225978 475494 226046
rect 474874 225922 474970 225978
rect 475026 225922 475094 225978
rect 475150 225922 475218 225978
rect 475274 225922 475342 225978
rect 475398 225922 475494 225978
rect 474874 208350 475494 225922
rect 474874 208294 474970 208350
rect 475026 208294 475094 208350
rect 475150 208294 475218 208350
rect 475274 208294 475342 208350
rect 475398 208294 475494 208350
rect 474874 208226 475494 208294
rect 474874 208170 474970 208226
rect 475026 208170 475094 208226
rect 475150 208170 475218 208226
rect 475274 208170 475342 208226
rect 475398 208170 475494 208226
rect 474874 208102 475494 208170
rect 474874 208046 474970 208102
rect 475026 208046 475094 208102
rect 475150 208046 475218 208102
rect 475274 208046 475342 208102
rect 475398 208046 475494 208102
rect 474874 207978 475494 208046
rect 474874 207922 474970 207978
rect 475026 207922 475094 207978
rect 475150 207922 475218 207978
rect 475274 207922 475342 207978
rect 475398 207922 475494 207978
rect 474874 190350 475494 207922
rect 474874 190294 474970 190350
rect 475026 190294 475094 190350
rect 475150 190294 475218 190350
rect 475274 190294 475342 190350
rect 475398 190294 475494 190350
rect 474874 190226 475494 190294
rect 474874 190170 474970 190226
rect 475026 190170 475094 190226
rect 475150 190170 475218 190226
rect 475274 190170 475342 190226
rect 475398 190170 475494 190226
rect 474874 190102 475494 190170
rect 474874 190046 474970 190102
rect 475026 190046 475094 190102
rect 475150 190046 475218 190102
rect 475274 190046 475342 190102
rect 475398 190046 475494 190102
rect 474874 189978 475494 190046
rect 474874 189922 474970 189978
rect 475026 189922 475094 189978
rect 475150 189922 475218 189978
rect 475274 189922 475342 189978
rect 475398 189922 475494 189978
rect 474874 172350 475494 189922
rect 474874 172294 474970 172350
rect 475026 172294 475094 172350
rect 475150 172294 475218 172350
rect 475274 172294 475342 172350
rect 475398 172294 475494 172350
rect 474874 172226 475494 172294
rect 474874 172170 474970 172226
rect 475026 172170 475094 172226
rect 475150 172170 475218 172226
rect 475274 172170 475342 172226
rect 475398 172170 475494 172226
rect 474874 172102 475494 172170
rect 474874 172046 474970 172102
rect 475026 172046 475094 172102
rect 475150 172046 475218 172102
rect 475274 172046 475342 172102
rect 475398 172046 475494 172102
rect 474874 171978 475494 172046
rect 474874 171922 474970 171978
rect 475026 171922 475094 171978
rect 475150 171922 475218 171978
rect 475274 171922 475342 171978
rect 475398 171922 475494 171978
rect 474874 154350 475494 171922
rect 474874 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 475494 154350
rect 474874 154226 475494 154294
rect 474874 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 475494 154226
rect 474874 154102 475494 154170
rect 474874 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 475494 154102
rect 474874 153978 475494 154046
rect 474874 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 475494 153978
rect 474874 136350 475494 153922
rect 474874 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 475494 136350
rect 474874 136226 475494 136294
rect 474874 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 475494 136226
rect 474874 136102 475494 136170
rect 474874 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 475494 136102
rect 474874 135978 475494 136046
rect 474874 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 475494 135978
rect 474874 118350 475494 135922
rect 474874 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 475494 118350
rect 474874 118226 475494 118294
rect 474874 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 475494 118226
rect 474874 118102 475494 118170
rect 474874 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 475494 118102
rect 474874 117978 475494 118046
rect 474874 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 475494 117978
rect 474874 100350 475494 117922
rect 474874 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 475494 100350
rect 474874 100226 475494 100294
rect 474874 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 475494 100226
rect 474874 100102 475494 100170
rect 474874 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 475494 100102
rect 474874 99978 475494 100046
rect 474874 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 475494 99978
rect 474874 82350 475494 99922
rect 474874 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 475494 82350
rect 474874 82226 475494 82294
rect 474874 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 475494 82226
rect 474874 82102 475494 82170
rect 474874 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 475494 82102
rect 474874 81978 475494 82046
rect 474874 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 475494 81978
rect 474874 64350 475494 81922
rect 474874 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 475494 64350
rect 474874 64226 475494 64294
rect 474874 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 475494 64226
rect 474874 64102 475494 64170
rect 474874 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 475494 64102
rect 474874 63978 475494 64046
rect 474874 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 475494 63978
rect 474874 46350 475494 63922
rect 474874 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 475494 46350
rect 474874 46226 475494 46294
rect 474874 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 475494 46226
rect 474874 46102 475494 46170
rect 474874 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 475494 46102
rect 474874 45978 475494 46046
rect 474874 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 475494 45978
rect 474874 28350 475494 45922
rect 474874 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 475494 28350
rect 474874 28226 475494 28294
rect 474874 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 475494 28226
rect 474874 28102 475494 28170
rect 474874 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 475494 28102
rect 474874 27978 475494 28046
rect 474874 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 475494 27978
rect 474874 10350 475494 27922
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 526350 489774 543922
rect 489154 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 489774 526350
rect 489154 526226 489774 526294
rect 489154 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 489774 526226
rect 489154 526102 489774 526170
rect 489154 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 489774 526102
rect 489154 525978 489774 526046
rect 489154 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 489774 525978
rect 489154 508350 489774 525922
rect 489154 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 489774 508350
rect 489154 508226 489774 508294
rect 489154 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 489774 508226
rect 489154 508102 489774 508170
rect 489154 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 489774 508102
rect 489154 507978 489774 508046
rect 489154 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 489774 507978
rect 489154 490350 489774 507922
rect 489154 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 489774 490350
rect 489154 490226 489774 490294
rect 489154 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 489774 490226
rect 489154 490102 489774 490170
rect 489154 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 489774 490102
rect 489154 489978 489774 490046
rect 489154 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 489774 489978
rect 489154 472350 489774 489922
rect 489154 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 489774 472350
rect 489154 472226 489774 472294
rect 489154 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 489774 472226
rect 489154 472102 489774 472170
rect 489154 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 489774 472102
rect 489154 471978 489774 472046
rect 489154 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 489774 471978
rect 489154 454350 489774 471922
rect 489154 454294 489250 454350
rect 489306 454294 489374 454350
rect 489430 454294 489498 454350
rect 489554 454294 489622 454350
rect 489678 454294 489774 454350
rect 489154 454226 489774 454294
rect 489154 454170 489250 454226
rect 489306 454170 489374 454226
rect 489430 454170 489498 454226
rect 489554 454170 489622 454226
rect 489678 454170 489774 454226
rect 489154 454102 489774 454170
rect 489154 454046 489250 454102
rect 489306 454046 489374 454102
rect 489430 454046 489498 454102
rect 489554 454046 489622 454102
rect 489678 454046 489774 454102
rect 489154 453978 489774 454046
rect 489154 453922 489250 453978
rect 489306 453922 489374 453978
rect 489430 453922 489498 453978
rect 489554 453922 489622 453978
rect 489678 453922 489774 453978
rect 489154 436350 489774 453922
rect 489154 436294 489250 436350
rect 489306 436294 489374 436350
rect 489430 436294 489498 436350
rect 489554 436294 489622 436350
rect 489678 436294 489774 436350
rect 489154 436226 489774 436294
rect 489154 436170 489250 436226
rect 489306 436170 489374 436226
rect 489430 436170 489498 436226
rect 489554 436170 489622 436226
rect 489678 436170 489774 436226
rect 489154 436102 489774 436170
rect 489154 436046 489250 436102
rect 489306 436046 489374 436102
rect 489430 436046 489498 436102
rect 489554 436046 489622 436102
rect 489678 436046 489774 436102
rect 489154 435978 489774 436046
rect 489154 435922 489250 435978
rect 489306 435922 489374 435978
rect 489430 435922 489498 435978
rect 489554 435922 489622 435978
rect 489678 435922 489774 435978
rect 489154 418350 489774 435922
rect 489154 418294 489250 418350
rect 489306 418294 489374 418350
rect 489430 418294 489498 418350
rect 489554 418294 489622 418350
rect 489678 418294 489774 418350
rect 489154 418226 489774 418294
rect 489154 418170 489250 418226
rect 489306 418170 489374 418226
rect 489430 418170 489498 418226
rect 489554 418170 489622 418226
rect 489678 418170 489774 418226
rect 489154 418102 489774 418170
rect 489154 418046 489250 418102
rect 489306 418046 489374 418102
rect 489430 418046 489498 418102
rect 489554 418046 489622 418102
rect 489678 418046 489774 418102
rect 489154 417978 489774 418046
rect 489154 417922 489250 417978
rect 489306 417922 489374 417978
rect 489430 417922 489498 417978
rect 489554 417922 489622 417978
rect 489678 417922 489774 417978
rect 489154 400350 489774 417922
rect 489154 400294 489250 400350
rect 489306 400294 489374 400350
rect 489430 400294 489498 400350
rect 489554 400294 489622 400350
rect 489678 400294 489774 400350
rect 489154 400226 489774 400294
rect 489154 400170 489250 400226
rect 489306 400170 489374 400226
rect 489430 400170 489498 400226
rect 489554 400170 489622 400226
rect 489678 400170 489774 400226
rect 489154 400102 489774 400170
rect 489154 400046 489250 400102
rect 489306 400046 489374 400102
rect 489430 400046 489498 400102
rect 489554 400046 489622 400102
rect 489678 400046 489774 400102
rect 489154 399978 489774 400046
rect 489154 399922 489250 399978
rect 489306 399922 489374 399978
rect 489430 399922 489498 399978
rect 489554 399922 489622 399978
rect 489678 399922 489774 399978
rect 489154 382350 489774 399922
rect 489154 382294 489250 382350
rect 489306 382294 489374 382350
rect 489430 382294 489498 382350
rect 489554 382294 489622 382350
rect 489678 382294 489774 382350
rect 489154 382226 489774 382294
rect 489154 382170 489250 382226
rect 489306 382170 489374 382226
rect 489430 382170 489498 382226
rect 489554 382170 489622 382226
rect 489678 382170 489774 382226
rect 489154 382102 489774 382170
rect 489154 382046 489250 382102
rect 489306 382046 489374 382102
rect 489430 382046 489498 382102
rect 489554 382046 489622 382102
rect 489678 382046 489774 382102
rect 489154 381978 489774 382046
rect 489154 381922 489250 381978
rect 489306 381922 489374 381978
rect 489430 381922 489498 381978
rect 489554 381922 489622 381978
rect 489678 381922 489774 381978
rect 489154 364350 489774 381922
rect 489154 364294 489250 364350
rect 489306 364294 489374 364350
rect 489430 364294 489498 364350
rect 489554 364294 489622 364350
rect 489678 364294 489774 364350
rect 489154 364226 489774 364294
rect 489154 364170 489250 364226
rect 489306 364170 489374 364226
rect 489430 364170 489498 364226
rect 489554 364170 489622 364226
rect 489678 364170 489774 364226
rect 489154 364102 489774 364170
rect 489154 364046 489250 364102
rect 489306 364046 489374 364102
rect 489430 364046 489498 364102
rect 489554 364046 489622 364102
rect 489678 364046 489774 364102
rect 489154 363978 489774 364046
rect 489154 363922 489250 363978
rect 489306 363922 489374 363978
rect 489430 363922 489498 363978
rect 489554 363922 489622 363978
rect 489678 363922 489774 363978
rect 489154 346350 489774 363922
rect 489154 346294 489250 346350
rect 489306 346294 489374 346350
rect 489430 346294 489498 346350
rect 489554 346294 489622 346350
rect 489678 346294 489774 346350
rect 489154 346226 489774 346294
rect 489154 346170 489250 346226
rect 489306 346170 489374 346226
rect 489430 346170 489498 346226
rect 489554 346170 489622 346226
rect 489678 346170 489774 346226
rect 489154 346102 489774 346170
rect 489154 346046 489250 346102
rect 489306 346046 489374 346102
rect 489430 346046 489498 346102
rect 489554 346046 489622 346102
rect 489678 346046 489774 346102
rect 489154 345978 489774 346046
rect 489154 345922 489250 345978
rect 489306 345922 489374 345978
rect 489430 345922 489498 345978
rect 489554 345922 489622 345978
rect 489678 345922 489774 345978
rect 489154 328350 489774 345922
rect 489154 328294 489250 328350
rect 489306 328294 489374 328350
rect 489430 328294 489498 328350
rect 489554 328294 489622 328350
rect 489678 328294 489774 328350
rect 489154 328226 489774 328294
rect 489154 328170 489250 328226
rect 489306 328170 489374 328226
rect 489430 328170 489498 328226
rect 489554 328170 489622 328226
rect 489678 328170 489774 328226
rect 489154 328102 489774 328170
rect 489154 328046 489250 328102
rect 489306 328046 489374 328102
rect 489430 328046 489498 328102
rect 489554 328046 489622 328102
rect 489678 328046 489774 328102
rect 489154 327978 489774 328046
rect 489154 327922 489250 327978
rect 489306 327922 489374 327978
rect 489430 327922 489498 327978
rect 489554 327922 489622 327978
rect 489678 327922 489774 327978
rect 489154 310350 489774 327922
rect 489154 310294 489250 310350
rect 489306 310294 489374 310350
rect 489430 310294 489498 310350
rect 489554 310294 489622 310350
rect 489678 310294 489774 310350
rect 489154 310226 489774 310294
rect 489154 310170 489250 310226
rect 489306 310170 489374 310226
rect 489430 310170 489498 310226
rect 489554 310170 489622 310226
rect 489678 310170 489774 310226
rect 489154 310102 489774 310170
rect 489154 310046 489250 310102
rect 489306 310046 489374 310102
rect 489430 310046 489498 310102
rect 489554 310046 489622 310102
rect 489678 310046 489774 310102
rect 489154 309978 489774 310046
rect 489154 309922 489250 309978
rect 489306 309922 489374 309978
rect 489430 309922 489498 309978
rect 489554 309922 489622 309978
rect 489678 309922 489774 309978
rect 489154 292350 489774 309922
rect 489154 292294 489250 292350
rect 489306 292294 489374 292350
rect 489430 292294 489498 292350
rect 489554 292294 489622 292350
rect 489678 292294 489774 292350
rect 489154 292226 489774 292294
rect 489154 292170 489250 292226
rect 489306 292170 489374 292226
rect 489430 292170 489498 292226
rect 489554 292170 489622 292226
rect 489678 292170 489774 292226
rect 489154 292102 489774 292170
rect 489154 292046 489250 292102
rect 489306 292046 489374 292102
rect 489430 292046 489498 292102
rect 489554 292046 489622 292102
rect 489678 292046 489774 292102
rect 489154 291978 489774 292046
rect 489154 291922 489250 291978
rect 489306 291922 489374 291978
rect 489430 291922 489498 291978
rect 489554 291922 489622 291978
rect 489678 291922 489774 291978
rect 489154 274350 489774 291922
rect 489154 274294 489250 274350
rect 489306 274294 489374 274350
rect 489430 274294 489498 274350
rect 489554 274294 489622 274350
rect 489678 274294 489774 274350
rect 489154 274226 489774 274294
rect 489154 274170 489250 274226
rect 489306 274170 489374 274226
rect 489430 274170 489498 274226
rect 489554 274170 489622 274226
rect 489678 274170 489774 274226
rect 489154 274102 489774 274170
rect 489154 274046 489250 274102
rect 489306 274046 489374 274102
rect 489430 274046 489498 274102
rect 489554 274046 489622 274102
rect 489678 274046 489774 274102
rect 489154 273978 489774 274046
rect 489154 273922 489250 273978
rect 489306 273922 489374 273978
rect 489430 273922 489498 273978
rect 489554 273922 489622 273978
rect 489678 273922 489774 273978
rect 489154 256350 489774 273922
rect 489154 256294 489250 256350
rect 489306 256294 489374 256350
rect 489430 256294 489498 256350
rect 489554 256294 489622 256350
rect 489678 256294 489774 256350
rect 489154 256226 489774 256294
rect 489154 256170 489250 256226
rect 489306 256170 489374 256226
rect 489430 256170 489498 256226
rect 489554 256170 489622 256226
rect 489678 256170 489774 256226
rect 489154 256102 489774 256170
rect 489154 256046 489250 256102
rect 489306 256046 489374 256102
rect 489430 256046 489498 256102
rect 489554 256046 489622 256102
rect 489678 256046 489774 256102
rect 489154 255978 489774 256046
rect 489154 255922 489250 255978
rect 489306 255922 489374 255978
rect 489430 255922 489498 255978
rect 489554 255922 489622 255978
rect 489678 255922 489774 255978
rect 489154 238350 489774 255922
rect 489154 238294 489250 238350
rect 489306 238294 489374 238350
rect 489430 238294 489498 238350
rect 489554 238294 489622 238350
rect 489678 238294 489774 238350
rect 489154 238226 489774 238294
rect 489154 238170 489250 238226
rect 489306 238170 489374 238226
rect 489430 238170 489498 238226
rect 489554 238170 489622 238226
rect 489678 238170 489774 238226
rect 489154 238102 489774 238170
rect 489154 238046 489250 238102
rect 489306 238046 489374 238102
rect 489430 238046 489498 238102
rect 489554 238046 489622 238102
rect 489678 238046 489774 238102
rect 489154 237978 489774 238046
rect 489154 237922 489250 237978
rect 489306 237922 489374 237978
rect 489430 237922 489498 237978
rect 489554 237922 489622 237978
rect 489678 237922 489774 237978
rect 489154 220350 489774 237922
rect 489154 220294 489250 220350
rect 489306 220294 489374 220350
rect 489430 220294 489498 220350
rect 489554 220294 489622 220350
rect 489678 220294 489774 220350
rect 489154 220226 489774 220294
rect 489154 220170 489250 220226
rect 489306 220170 489374 220226
rect 489430 220170 489498 220226
rect 489554 220170 489622 220226
rect 489678 220170 489774 220226
rect 489154 220102 489774 220170
rect 489154 220046 489250 220102
rect 489306 220046 489374 220102
rect 489430 220046 489498 220102
rect 489554 220046 489622 220102
rect 489678 220046 489774 220102
rect 489154 219978 489774 220046
rect 489154 219922 489250 219978
rect 489306 219922 489374 219978
rect 489430 219922 489498 219978
rect 489554 219922 489622 219978
rect 489678 219922 489774 219978
rect 489154 202350 489774 219922
rect 489154 202294 489250 202350
rect 489306 202294 489374 202350
rect 489430 202294 489498 202350
rect 489554 202294 489622 202350
rect 489678 202294 489774 202350
rect 489154 202226 489774 202294
rect 489154 202170 489250 202226
rect 489306 202170 489374 202226
rect 489430 202170 489498 202226
rect 489554 202170 489622 202226
rect 489678 202170 489774 202226
rect 489154 202102 489774 202170
rect 489154 202046 489250 202102
rect 489306 202046 489374 202102
rect 489430 202046 489498 202102
rect 489554 202046 489622 202102
rect 489678 202046 489774 202102
rect 489154 201978 489774 202046
rect 489154 201922 489250 201978
rect 489306 201922 489374 201978
rect 489430 201922 489498 201978
rect 489554 201922 489622 201978
rect 489678 201922 489774 201978
rect 489154 184350 489774 201922
rect 489154 184294 489250 184350
rect 489306 184294 489374 184350
rect 489430 184294 489498 184350
rect 489554 184294 489622 184350
rect 489678 184294 489774 184350
rect 489154 184226 489774 184294
rect 489154 184170 489250 184226
rect 489306 184170 489374 184226
rect 489430 184170 489498 184226
rect 489554 184170 489622 184226
rect 489678 184170 489774 184226
rect 489154 184102 489774 184170
rect 489154 184046 489250 184102
rect 489306 184046 489374 184102
rect 489430 184046 489498 184102
rect 489554 184046 489622 184102
rect 489678 184046 489774 184102
rect 489154 183978 489774 184046
rect 489154 183922 489250 183978
rect 489306 183922 489374 183978
rect 489430 183922 489498 183978
rect 489554 183922 489622 183978
rect 489678 183922 489774 183978
rect 489154 166350 489774 183922
rect 489154 166294 489250 166350
rect 489306 166294 489374 166350
rect 489430 166294 489498 166350
rect 489554 166294 489622 166350
rect 489678 166294 489774 166350
rect 489154 166226 489774 166294
rect 489154 166170 489250 166226
rect 489306 166170 489374 166226
rect 489430 166170 489498 166226
rect 489554 166170 489622 166226
rect 489678 166170 489774 166226
rect 489154 166102 489774 166170
rect 489154 166046 489250 166102
rect 489306 166046 489374 166102
rect 489430 166046 489498 166102
rect 489554 166046 489622 166102
rect 489678 166046 489774 166102
rect 489154 165978 489774 166046
rect 489154 165922 489250 165978
rect 489306 165922 489374 165978
rect 489430 165922 489498 165978
rect 489554 165922 489622 165978
rect 489678 165922 489774 165978
rect 489154 148350 489774 165922
rect 489154 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 489774 148350
rect 489154 148226 489774 148294
rect 489154 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 489774 148226
rect 489154 148102 489774 148170
rect 489154 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 489774 148102
rect 489154 147978 489774 148046
rect 489154 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 489774 147978
rect 489154 130350 489774 147922
rect 489154 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 489774 130350
rect 489154 130226 489774 130294
rect 489154 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 489774 130226
rect 489154 130102 489774 130170
rect 489154 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 489774 130102
rect 489154 129978 489774 130046
rect 489154 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 489774 129978
rect 489154 112350 489774 129922
rect 489154 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 489774 112350
rect 489154 112226 489774 112294
rect 489154 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 489774 112226
rect 489154 112102 489774 112170
rect 489154 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 489774 112102
rect 489154 111978 489774 112046
rect 489154 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 489774 111978
rect 489154 94350 489774 111922
rect 489154 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 489774 94350
rect 489154 94226 489774 94294
rect 489154 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 489774 94226
rect 489154 94102 489774 94170
rect 489154 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 489774 94102
rect 489154 93978 489774 94046
rect 489154 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 489774 93978
rect 489154 76350 489774 93922
rect 489154 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 489774 76350
rect 489154 76226 489774 76294
rect 489154 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 489774 76226
rect 489154 76102 489774 76170
rect 489154 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 489774 76102
rect 489154 75978 489774 76046
rect 489154 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 489774 75978
rect 489154 58350 489774 75922
rect 489154 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 489774 58350
rect 489154 58226 489774 58294
rect 489154 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 489774 58226
rect 489154 58102 489774 58170
rect 489154 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 489774 58102
rect 489154 57978 489774 58046
rect 489154 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 489774 57978
rect 489154 40350 489774 57922
rect 489154 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 489774 40350
rect 489154 40226 489774 40294
rect 489154 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 489774 40226
rect 489154 40102 489774 40170
rect 489154 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 489774 40102
rect 489154 39978 489774 40046
rect 489154 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 489774 39978
rect 489154 22350 489774 39922
rect 489154 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 489774 22350
rect 489154 22226 489774 22294
rect 489154 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 489774 22226
rect 489154 22102 489774 22170
rect 489154 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 489774 22102
rect 489154 21978 489774 22046
rect 489154 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 489774 21978
rect 489154 4350 489774 21922
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 514350 493494 531922
rect 492874 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 493494 514350
rect 492874 514226 493494 514294
rect 492874 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 493494 514226
rect 492874 514102 493494 514170
rect 492874 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 493494 514102
rect 492874 513978 493494 514046
rect 492874 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 493494 513978
rect 492874 496350 493494 513922
rect 492874 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 493494 496350
rect 492874 496226 493494 496294
rect 492874 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 493494 496226
rect 492874 496102 493494 496170
rect 492874 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 493494 496102
rect 492874 495978 493494 496046
rect 492874 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 493494 495978
rect 492874 478350 493494 495922
rect 492874 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 493494 478350
rect 492874 478226 493494 478294
rect 492874 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 493494 478226
rect 492874 478102 493494 478170
rect 492874 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 493494 478102
rect 492874 477978 493494 478046
rect 492874 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 493494 477978
rect 492874 460350 493494 477922
rect 492874 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 493494 460350
rect 492874 460226 493494 460294
rect 492874 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 493494 460226
rect 492874 460102 493494 460170
rect 492874 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 493494 460102
rect 492874 459978 493494 460046
rect 492874 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 493494 459978
rect 492874 442350 493494 459922
rect 492874 442294 492970 442350
rect 493026 442294 493094 442350
rect 493150 442294 493218 442350
rect 493274 442294 493342 442350
rect 493398 442294 493494 442350
rect 492874 442226 493494 442294
rect 492874 442170 492970 442226
rect 493026 442170 493094 442226
rect 493150 442170 493218 442226
rect 493274 442170 493342 442226
rect 493398 442170 493494 442226
rect 492874 442102 493494 442170
rect 492874 442046 492970 442102
rect 493026 442046 493094 442102
rect 493150 442046 493218 442102
rect 493274 442046 493342 442102
rect 493398 442046 493494 442102
rect 492874 441978 493494 442046
rect 492874 441922 492970 441978
rect 493026 441922 493094 441978
rect 493150 441922 493218 441978
rect 493274 441922 493342 441978
rect 493398 441922 493494 441978
rect 492874 424350 493494 441922
rect 492874 424294 492970 424350
rect 493026 424294 493094 424350
rect 493150 424294 493218 424350
rect 493274 424294 493342 424350
rect 493398 424294 493494 424350
rect 492874 424226 493494 424294
rect 492874 424170 492970 424226
rect 493026 424170 493094 424226
rect 493150 424170 493218 424226
rect 493274 424170 493342 424226
rect 493398 424170 493494 424226
rect 492874 424102 493494 424170
rect 492874 424046 492970 424102
rect 493026 424046 493094 424102
rect 493150 424046 493218 424102
rect 493274 424046 493342 424102
rect 493398 424046 493494 424102
rect 492874 423978 493494 424046
rect 492874 423922 492970 423978
rect 493026 423922 493094 423978
rect 493150 423922 493218 423978
rect 493274 423922 493342 423978
rect 493398 423922 493494 423978
rect 492874 406350 493494 423922
rect 492874 406294 492970 406350
rect 493026 406294 493094 406350
rect 493150 406294 493218 406350
rect 493274 406294 493342 406350
rect 493398 406294 493494 406350
rect 492874 406226 493494 406294
rect 492874 406170 492970 406226
rect 493026 406170 493094 406226
rect 493150 406170 493218 406226
rect 493274 406170 493342 406226
rect 493398 406170 493494 406226
rect 492874 406102 493494 406170
rect 492874 406046 492970 406102
rect 493026 406046 493094 406102
rect 493150 406046 493218 406102
rect 493274 406046 493342 406102
rect 493398 406046 493494 406102
rect 492874 405978 493494 406046
rect 492874 405922 492970 405978
rect 493026 405922 493094 405978
rect 493150 405922 493218 405978
rect 493274 405922 493342 405978
rect 493398 405922 493494 405978
rect 492874 388350 493494 405922
rect 492874 388294 492970 388350
rect 493026 388294 493094 388350
rect 493150 388294 493218 388350
rect 493274 388294 493342 388350
rect 493398 388294 493494 388350
rect 492874 388226 493494 388294
rect 492874 388170 492970 388226
rect 493026 388170 493094 388226
rect 493150 388170 493218 388226
rect 493274 388170 493342 388226
rect 493398 388170 493494 388226
rect 492874 388102 493494 388170
rect 492874 388046 492970 388102
rect 493026 388046 493094 388102
rect 493150 388046 493218 388102
rect 493274 388046 493342 388102
rect 493398 388046 493494 388102
rect 492874 387978 493494 388046
rect 492874 387922 492970 387978
rect 493026 387922 493094 387978
rect 493150 387922 493218 387978
rect 493274 387922 493342 387978
rect 493398 387922 493494 387978
rect 492874 370350 493494 387922
rect 492874 370294 492970 370350
rect 493026 370294 493094 370350
rect 493150 370294 493218 370350
rect 493274 370294 493342 370350
rect 493398 370294 493494 370350
rect 492874 370226 493494 370294
rect 492874 370170 492970 370226
rect 493026 370170 493094 370226
rect 493150 370170 493218 370226
rect 493274 370170 493342 370226
rect 493398 370170 493494 370226
rect 492874 370102 493494 370170
rect 492874 370046 492970 370102
rect 493026 370046 493094 370102
rect 493150 370046 493218 370102
rect 493274 370046 493342 370102
rect 493398 370046 493494 370102
rect 492874 369978 493494 370046
rect 492874 369922 492970 369978
rect 493026 369922 493094 369978
rect 493150 369922 493218 369978
rect 493274 369922 493342 369978
rect 493398 369922 493494 369978
rect 492874 352350 493494 369922
rect 492874 352294 492970 352350
rect 493026 352294 493094 352350
rect 493150 352294 493218 352350
rect 493274 352294 493342 352350
rect 493398 352294 493494 352350
rect 492874 352226 493494 352294
rect 492874 352170 492970 352226
rect 493026 352170 493094 352226
rect 493150 352170 493218 352226
rect 493274 352170 493342 352226
rect 493398 352170 493494 352226
rect 492874 352102 493494 352170
rect 492874 352046 492970 352102
rect 493026 352046 493094 352102
rect 493150 352046 493218 352102
rect 493274 352046 493342 352102
rect 493398 352046 493494 352102
rect 492874 351978 493494 352046
rect 492874 351922 492970 351978
rect 493026 351922 493094 351978
rect 493150 351922 493218 351978
rect 493274 351922 493342 351978
rect 493398 351922 493494 351978
rect 492874 334350 493494 351922
rect 492874 334294 492970 334350
rect 493026 334294 493094 334350
rect 493150 334294 493218 334350
rect 493274 334294 493342 334350
rect 493398 334294 493494 334350
rect 492874 334226 493494 334294
rect 492874 334170 492970 334226
rect 493026 334170 493094 334226
rect 493150 334170 493218 334226
rect 493274 334170 493342 334226
rect 493398 334170 493494 334226
rect 492874 334102 493494 334170
rect 492874 334046 492970 334102
rect 493026 334046 493094 334102
rect 493150 334046 493218 334102
rect 493274 334046 493342 334102
rect 493398 334046 493494 334102
rect 492874 333978 493494 334046
rect 492874 333922 492970 333978
rect 493026 333922 493094 333978
rect 493150 333922 493218 333978
rect 493274 333922 493342 333978
rect 493398 333922 493494 333978
rect 492874 316350 493494 333922
rect 492874 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 493494 316350
rect 492874 316226 493494 316294
rect 492874 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 493494 316226
rect 492874 316102 493494 316170
rect 492874 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 493494 316102
rect 492874 315978 493494 316046
rect 492874 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 493494 315978
rect 492874 298350 493494 315922
rect 492874 298294 492970 298350
rect 493026 298294 493094 298350
rect 493150 298294 493218 298350
rect 493274 298294 493342 298350
rect 493398 298294 493494 298350
rect 492874 298226 493494 298294
rect 492874 298170 492970 298226
rect 493026 298170 493094 298226
rect 493150 298170 493218 298226
rect 493274 298170 493342 298226
rect 493398 298170 493494 298226
rect 492874 298102 493494 298170
rect 492874 298046 492970 298102
rect 493026 298046 493094 298102
rect 493150 298046 493218 298102
rect 493274 298046 493342 298102
rect 493398 298046 493494 298102
rect 492874 297978 493494 298046
rect 492874 297922 492970 297978
rect 493026 297922 493094 297978
rect 493150 297922 493218 297978
rect 493274 297922 493342 297978
rect 493398 297922 493494 297978
rect 492874 280350 493494 297922
rect 492874 280294 492970 280350
rect 493026 280294 493094 280350
rect 493150 280294 493218 280350
rect 493274 280294 493342 280350
rect 493398 280294 493494 280350
rect 492874 280226 493494 280294
rect 492874 280170 492970 280226
rect 493026 280170 493094 280226
rect 493150 280170 493218 280226
rect 493274 280170 493342 280226
rect 493398 280170 493494 280226
rect 492874 280102 493494 280170
rect 492874 280046 492970 280102
rect 493026 280046 493094 280102
rect 493150 280046 493218 280102
rect 493274 280046 493342 280102
rect 493398 280046 493494 280102
rect 492874 279978 493494 280046
rect 492874 279922 492970 279978
rect 493026 279922 493094 279978
rect 493150 279922 493218 279978
rect 493274 279922 493342 279978
rect 493398 279922 493494 279978
rect 492874 262350 493494 279922
rect 492874 262294 492970 262350
rect 493026 262294 493094 262350
rect 493150 262294 493218 262350
rect 493274 262294 493342 262350
rect 493398 262294 493494 262350
rect 492874 262226 493494 262294
rect 492874 262170 492970 262226
rect 493026 262170 493094 262226
rect 493150 262170 493218 262226
rect 493274 262170 493342 262226
rect 493398 262170 493494 262226
rect 492874 262102 493494 262170
rect 492874 262046 492970 262102
rect 493026 262046 493094 262102
rect 493150 262046 493218 262102
rect 493274 262046 493342 262102
rect 493398 262046 493494 262102
rect 492874 261978 493494 262046
rect 492874 261922 492970 261978
rect 493026 261922 493094 261978
rect 493150 261922 493218 261978
rect 493274 261922 493342 261978
rect 493398 261922 493494 261978
rect 492874 244350 493494 261922
rect 492874 244294 492970 244350
rect 493026 244294 493094 244350
rect 493150 244294 493218 244350
rect 493274 244294 493342 244350
rect 493398 244294 493494 244350
rect 492874 244226 493494 244294
rect 492874 244170 492970 244226
rect 493026 244170 493094 244226
rect 493150 244170 493218 244226
rect 493274 244170 493342 244226
rect 493398 244170 493494 244226
rect 492874 244102 493494 244170
rect 492874 244046 492970 244102
rect 493026 244046 493094 244102
rect 493150 244046 493218 244102
rect 493274 244046 493342 244102
rect 493398 244046 493494 244102
rect 492874 243978 493494 244046
rect 492874 243922 492970 243978
rect 493026 243922 493094 243978
rect 493150 243922 493218 243978
rect 493274 243922 493342 243978
rect 493398 243922 493494 243978
rect 492874 226350 493494 243922
rect 492874 226294 492970 226350
rect 493026 226294 493094 226350
rect 493150 226294 493218 226350
rect 493274 226294 493342 226350
rect 493398 226294 493494 226350
rect 492874 226226 493494 226294
rect 492874 226170 492970 226226
rect 493026 226170 493094 226226
rect 493150 226170 493218 226226
rect 493274 226170 493342 226226
rect 493398 226170 493494 226226
rect 492874 226102 493494 226170
rect 492874 226046 492970 226102
rect 493026 226046 493094 226102
rect 493150 226046 493218 226102
rect 493274 226046 493342 226102
rect 493398 226046 493494 226102
rect 492874 225978 493494 226046
rect 492874 225922 492970 225978
rect 493026 225922 493094 225978
rect 493150 225922 493218 225978
rect 493274 225922 493342 225978
rect 493398 225922 493494 225978
rect 492874 208350 493494 225922
rect 492874 208294 492970 208350
rect 493026 208294 493094 208350
rect 493150 208294 493218 208350
rect 493274 208294 493342 208350
rect 493398 208294 493494 208350
rect 492874 208226 493494 208294
rect 492874 208170 492970 208226
rect 493026 208170 493094 208226
rect 493150 208170 493218 208226
rect 493274 208170 493342 208226
rect 493398 208170 493494 208226
rect 492874 208102 493494 208170
rect 492874 208046 492970 208102
rect 493026 208046 493094 208102
rect 493150 208046 493218 208102
rect 493274 208046 493342 208102
rect 493398 208046 493494 208102
rect 492874 207978 493494 208046
rect 492874 207922 492970 207978
rect 493026 207922 493094 207978
rect 493150 207922 493218 207978
rect 493274 207922 493342 207978
rect 493398 207922 493494 207978
rect 492874 190350 493494 207922
rect 492874 190294 492970 190350
rect 493026 190294 493094 190350
rect 493150 190294 493218 190350
rect 493274 190294 493342 190350
rect 493398 190294 493494 190350
rect 492874 190226 493494 190294
rect 492874 190170 492970 190226
rect 493026 190170 493094 190226
rect 493150 190170 493218 190226
rect 493274 190170 493342 190226
rect 493398 190170 493494 190226
rect 492874 190102 493494 190170
rect 492874 190046 492970 190102
rect 493026 190046 493094 190102
rect 493150 190046 493218 190102
rect 493274 190046 493342 190102
rect 493398 190046 493494 190102
rect 492874 189978 493494 190046
rect 492874 189922 492970 189978
rect 493026 189922 493094 189978
rect 493150 189922 493218 189978
rect 493274 189922 493342 189978
rect 493398 189922 493494 189978
rect 492874 172350 493494 189922
rect 492874 172294 492970 172350
rect 493026 172294 493094 172350
rect 493150 172294 493218 172350
rect 493274 172294 493342 172350
rect 493398 172294 493494 172350
rect 492874 172226 493494 172294
rect 492874 172170 492970 172226
rect 493026 172170 493094 172226
rect 493150 172170 493218 172226
rect 493274 172170 493342 172226
rect 493398 172170 493494 172226
rect 492874 172102 493494 172170
rect 492874 172046 492970 172102
rect 493026 172046 493094 172102
rect 493150 172046 493218 172102
rect 493274 172046 493342 172102
rect 493398 172046 493494 172102
rect 492874 171978 493494 172046
rect 492874 171922 492970 171978
rect 493026 171922 493094 171978
rect 493150 171922 493218 171978
rect 493274 171922 493342 171978
rect 493398 171922 493494 171978
rect 492874 154350 493494 171922
rect 492874 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 493494 154350
rect 492874 154226 493494 154294
rect 492874 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 493494 154226
rect 492874 154102 493494 154170
rect 492874 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 493494 154102
rect 492874 153978 493494 154046
rect 492874 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 493494 153978
rect 492874 136350 493494 153922
rect 492874 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 493494 136350
rect 492874 136226 493494 136294
rect 492874 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 493494 136226
rect 492874 136102 493494 136170
rect 492874 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 493494 136102
rect 492874 135978 493494 136046
rect 492874 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 493494 135978
rect 492874 118350 493494 135922
rect 492874 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 493494 118350
rect 492874 118226 493494 118294
rect 492874 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 493494 118226
rect 492874 118102 493494 118170
rect 492874 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 493494 118102
rect 492874 117978 493494 118046
rect 492874 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 493494 117978
rect 492874 100350 493494 117922
rect 492874 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 493494 100350
rect 492874 100226 493494 100294
rect 492874 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 493494 100226
rect 492874 100102 493494 100170
rect 492874 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 493494 100102
rect 492874 99978 493494 100046
rect 492874 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 493494 99978
rect 492874 82350 493494 99922
rect 492874 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 493494 82350
rect 492874 82226 493494 82294
rect 492874 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 493494 82226
rect 492874 82102 493494 82170
rect 492874 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 493494 82102
rect 492874 81978 493494 82046
rect 492874 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 493494 81978
rect 492874 64350 493494 81922
rect 492874 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 493494 64350
rect 492874 64226 493494 64294
rect 492874 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 493494 64226
rect 492874 64102 493494 64170
rect 492874 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 493494 64102
rect 492874 63978 493494 64046
rect 492874 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 493494 63978
rect 492874 46350 493494 63922
rect 492874 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 493494 46350
rect 492874 46226 493494 46294
rect 492874 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 493494 46226
rect 492874 46102 493494 46170
rect 492874 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 493494 46102
rect 492874 45978 493494 46046
rect 492874 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 493494 45978
rect 492874 28350 493494 45922
rect 492874 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 493494 28350
rect 492874 28226 493494 28294
rect 492874 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 493494 28226
rect 492874 28102 493494 28170
rect 492874 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 493494 28102
rect 492874 27978 493494 28046
rect 492874 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 493494 27978
rect 492874 10350 493494 27922
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 526350 507774 543922
rect 507154 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 507774 526350
rect 507154 526226 507774 526294
rect 507154 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 507774 526226
rect 507154 526102 507774 526170
rect 507154 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 507774 526102
rect 507154 525978 507774 526046
rect 507154 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 507774 525978
rect 507154 508350 507774 525922
rect 507154 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 507774 508350
rect 507154 508226 507774 508294
rect 507154 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 507774 508226
rect 507154 508102 507774 508170
rect 507154 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 507774 508102
rect 507154 507978 507774 508046
rect 507154 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 507774 507978
rect 507154 490350 507774 507922
rect 507154 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 507774 490350
rect 507154 490226 507774 490294
rect 507154 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 507774 490226
rect 507154 490102 507774 490170
rect 507154 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 507774 490102
rect 507154 489978 507774 490046
rect 507154 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 507774 489978
rect 507154 472350 507774 489922
rect 507154 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 507774 472350
rect 507154 472226 507774 472294
rect 507154 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 507774 472226
rect 507154 472102 507774 472170
rect 507154 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 507774 472102
rect 507154 471978 507774 472046
rect 507154 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 507774 471978
rect 507154 454350 507774 471922
rect 507154 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 507774 454350
rect 507154 454226 507774 454294
rect 507154 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 507774 454226
rect 507154 454102 507774 454170
rect 507154 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 507774 454102
rect 507154 453978 507774 454046
rect 507154 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 507774 453978
rect 507154 436350 507774 453922
rect 507154 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 507774 436350
rect 507154 436226 507774 436294
rect 507154 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 507774 436226
rect 507154 436102 507774 436170
rect 507154 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 507774 436102
rect 507154 435978 507774 436046
rect 507154 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 507774 435978
rect 507154 418350 507774 435922
rect 507154 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 507774 418350
rect 507154 418226 507774 418294
rect 507154 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 507774 418226
rect 507154 418102 507774 418170
rect 507154 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 507774 418102
rect 507154 417978 507774 418046
rect 507154 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 507774 417978
rect 507154 400350 507774 417922
rect 507154 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 507774 400350
rect 507154 400226 507774 400294
rect 507154 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 507774 400226
rect 507154 400102 507774 400170
rect 507154 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 507774 400102
rect 507154 399978 507774 400046
rect 507154 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 507774 399978
rect 507154 382350 507774 399922
rect 507154 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 507774 382350
rect 507154 382226 507774 382294
rect 507154 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 507774 382226
rect 507154 382102 507774 382170
rect 507154 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 507774 382102
rect 507154 381978 507774 382046
rect 507154 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 507774 381978
rect 507154 364350 507774 381922
rect 507154 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 507774 364350
rect 507154 364226 507774 364294
rect 507154 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 507774 364226
rect 507154 364102 507774 364170
rect 507154 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 507774 364102
rect 507154 363978 507774 364046
rect 507154 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 507774 363978
rect 507154 346350 507774 363922
rect 507154 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 507774 346350
rect 507154 346226 507774 346294
rect 507154 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 507774 346226
rect 507154 346102 507774 346170
rect 507154 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 507774 346102
rect 507154 345978 507774 346046
rect 507154 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 507774 345978
rect 507154 328350 507774 345922
rect 507154 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 507774 328350
rect 507154 328226 507774 328294
rect 507154 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 507774 328226
rect 507154 328102 507774 328170
rect 507154 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 507774 328102
rect 507154 327978 507774 328046
rect 507154 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 507774 327978
rect 507154 310350 507774 327922
rect 507154 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 507774 310350
rect 507154 310226 507774 310294
rect 507154 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 507774 310226
rect 507154 310102 507774 310170
rect 507154 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 507774 310102
rect 507154 309978 507774 310046
rect 507154 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 507774 309978
rect 507154 292350 507774 309922
rect 507154 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 507774 292350
rect 507154 292226 507774 292294
rect 507154 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 507774 292226
rect 507154 292102 507774 292170
rect 507154 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 507774 292102
rect 507154 291978 507774 292046
rect 507154 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 507774 291978
rect 507154 274350 507774 291922
rect 507154 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 507774 274350
rect 507154 274226 507774 274294
rect 507154 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 507774 274226
rect 507154 274102 507774 274170
rect 507154 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 507774 274102
rect 507154 273978 507774 274046
rect 507154 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 507774 273978
rect 507154 256350 507774 273922
rect 507154 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 507774 256350
rect 507154 256226 507774 256294
rect 507154 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 507774 256226
rect 507154 256102 507774 256170
rect 507154 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 507774 256102
rect 507154 255978 507774 256046
rect 507154 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 507774 255978
rect 507154 238350 507774 255922
rect 507154 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 507774 238350
rect 507154 238226 507774 238294
rect 507154 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 507774 238226
rect 507154 238102 507774 238170
rect 507154 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 507774 238102
rect 507154 237978 507774 238046
rect 507154 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 507774 237978
rect 507154 220350 507774 237922
rect 507154 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 507774 220350
rect 507154 220226 507774 220294
rect 507154 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 507774 220226
rect 507154 220102 507774 220170
rect 507154 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 507774 220102
rect 507154 219978 507774 220046
rect 507154 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 507774 219978
rect 507154 202350 507774 219922
rect 507154 202294 507250 202350
rect 507306 202294 507374 202350
rect 507430 202294 507498 202350
rect 507554 202294 507622 202350
rect 507678 202294 507774 202350
rect 507154 202226 507774 202294
rect 507154 202170 507250 202226
rect 507306 202170 507374 202226
rect 507430 202170 507498 202226
rect 507554 202170 507622 202226
rect 507678 202170 507774 202226
rect 507154 202102 507774 202170
rect 507154 202046 507250 202102
rect 507306 202046 507374 202102
rect 507430 202046 507498 202102
rect 507554 202046 507622 202102
rect 507678 202046 507774 202102
rect 507154 201978 507774 202046
rect 507154 201922 507250 201978
rect 507306 201922 507374 201978
rect 507430 201922 507498 201978
rect 507554 201922 507622 201978
rect 507678 201922 507774 201978
rect 507154 184350 507774 201922
rect 507154 184294 507250 184350
rect 507306 184294 507374 184350
rect 507430 184294 507498 184350
rect 507554 184294 507622 184350
rect 507678 184294 507774 184350
rect 507154 184226 507774 184294
rect 507154 184170 507250 184226
rect 507306 184170 507374 184226
rect 507430 184170 507498 184226
rect 507554 184170 507622 184226
rect 507678 184170 507774 184226
rect 507154 184102 507774 184170
rect 507154 184046 507250 184102
rect 507306 184046 507374 184102
rect 507430 184046 507498 184102
rect 507554 184046 507622 184102
rect 507678 184046 507774 184102
rect 507154 183978 507774 184046
rect 507154 183922 507250 183978
rect 507306 183922 507374 183978
rect 507430 183922 507498 183978
rect 507554 183922 507622 183978
rect 507678 183922 507774 183978
rect 507154 166350 507774 183922
rect 507154 166294 507250 166350
rect 507306 166294 507374 166350
rect 507430 166294 507498 166350
rect 507554 166294 507622 166350
rect 507678 166294 507774 166350
rect 507154 166226 507774 166294
rect 507154 166170 507250 166226
rect 507306 166170 507374 166226
rect 507430 166170 507498 166226
rect 507554 166170 507622 166226
rect 507678 166170 507774 166226
rect 507154 166102 507774 166170
rect 507154 166046 507250 166102
rect 507306 166046 507374 166102
rect 507430 166046 507498 166102
rect 507554 166046 507622 166102
rect 507678 166046 507774 166102
rect 507154 165978 507774 166046
rect 507154 165922 507250 165978
rect 507306 165922 507374 165978
rect 507430 165922 507498 165978
rect 507554 165922 507622 165978
rect 507678 165922 507774 165978
rect 507154 148350 507774 165922
rect 507154 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 507774 148350
rect 507154 148226 507774 148294
rect 507154 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 507774 148226
rect 507154 148102 507774 148170
rect 507154 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 507774 148102
rect 507154 147978 507774 148046
rect 507154 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 507774 147978
rect 507154 130350 507774 147922
rect 507154 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 507774 130350
rect 507154 130226 507774 130294
rect 507154 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 507774 130226
rect 507154 130102 507774 130170
rect 507154 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 507774 130102
rect 507154 129978 507774 130046
rect 507154 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 507774 129978
rect 507154 112350 507774 129922
rect 507154 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 507774 112350
rect 507154 112226 507774 112294
rect 507154 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 507774 112226
rect 507154 112102 507774 112170
rect 507154 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 507774 112102
rect 507154 111978 507774 112046
rect 507154 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 507774 111978
rect 507154 94350 507774 111922
rect 507154 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 507774 94350
rect 507154 94226 507774 94294
rect 507154 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 507774 94226
rect 507154 94102 507774 94170
rect 507154 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 507774 94102
rect 507154 93978 507774 94046
rect 507154 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 507774 93978
rect 507154 76350 507774 93922
rect 507154 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 507774 76350
rect 507154 76226 507774 76294
rect 507154 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 507774 76226
rect 507154 76102 507774 76170
rect 507154 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 507774 76102
rect 507154 75978 507774 76046
rect 507154 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 507774 75978
rect 507154 58350 507774 75922
rect 507154 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 507774 58350
rect 507154 58226 507774 58294
rect 507154 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 507774 58226
rect 507154 58102 507774 58170
rect 507154 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 507774 58102
rect 507154 57978 507774 58046
rect 507154 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 507774 57978
rect 507154 40350 507774 57922
rect 507154 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 507774 40350
rect 507154 40226 507774 40294
rect 507154 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 507774 40226
rect 507154 40102 507774 40170
rect 507154 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 507774 40102
rect 507154 39978 507774 40046
rect 507154 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 507774 39978
rect 507154 22350 507774 39922
rect 507154 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 507774 22350
rect 507154 22226 507774 22294
rect 507154 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 507774 22226
rect 507154 22102 507774 22170
rect 507154 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 507774 22102
rect 507154 21978 507774 22046
rect 507154 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 507774 21978
rect 507154 4350 507774 21922
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 514350 511494 531922
rect 510874 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 511494 514350
rect 510874 514226 511494 514294
rect 510874 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 511494 514226
rect 510874 514102 511494 514170
rect 510874 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 511494 514102
rect 510874 513978 511494 514046
rect 510874 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 511494 513978
rect 510874 496350 511494 513922
rect 510874 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 511494 496350
rect 510874 496226 511494 496294
rect 510874 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 511494 496226
rect 510874 496102 511494 496170
rect 510874 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 511494 496102
rect 510874 495978 511494 496046
rect 510874 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 511494 495978
rect 510874 478350 511494 495922
rect 510874 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 511494 478350
rect 510874 478226 511494 478294
rect 510874 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 511494 478226
rect 510874 478102 511494 478170
rect 510874 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 511494 478102
rect 510874 477978 511494 478046
rect 510874 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 511494 477978
rect 510874 460350 511494 477922
rect 510874 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 511494 460350
rect 510874 460226 511494 460294
rect 510874 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 511494 460226
rect 510874 460102 511494 460170
rect 510874 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 511494 460102
rect 510874 459978 511494 460046
rect 510874 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 511494 459978
rect 510874 442350 511494 459922
rect 510874 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 511494 442350
rect 510874 442226 511494 442294
rect 510874 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 511494 442226
rect 510874 442102 511494 442170
rect 510874 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 511494 442102
rect 510874 441978 511494 442046
rect 510874 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 511494 441978
rect 510874 424350 511494 441922
rect 510874 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 511494 424350
rect 510874 424226 511494 424294
rect 510874 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 511494 424226
rect 510874 424102 511494 424170
rect 510874 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 511494 424102
rect 510874 423978 511494 424046
rect 510874 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 511494 423978
rect 510874 406350 511494 423922
rect 510874 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 511494 406350
rect 510874 406226 511494 406294
rect 510874 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 511494 406226
rect 510874 406102 511494 406170
rect 510874 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 511494 406102
rect 510874 405978 511494 406046
rect 510874 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 511494 405978
rect 510874 388350 511494 405922
rect 510874 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 511494 388350
rect 510874 388226 511494 388294
rect 510874 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 511494 388226
rect 510874 388102 511494 388170
rect 510874 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 511494 388102
rect 510874 387978 511494 388046
rect 510874 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 511494 387978
rect 510874 370350 511494 387922
rect 510874 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 511494 370350
rect 510874 370226 511494 370294
rect 510874 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 511494 370226
rect 510874 370102 511494 370170
rect 510874 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 511494 370102
rect 510874 369978 511494 370046
rect 510874 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 511494 369978
rect 510874 352350 511494 369922
rect 510874 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 511494 352350
rect 510874 352226 511494 352294
rect 510874 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 511494 352226
rect 510874 352102 511494 352170
rect 510874 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 511494 352102
rect 510874 351978 511494 352046
rect 510874 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 511494 351978
rect 510874 334350 511494 351922
rect 510874 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 511494 334350
rect 510874 334226 511494 334294
rect 510874 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 511494 334226
rect 510874 334102 511494 334170
rect 510874 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 511494 334102
rect 510874 333978 511494 334046
rect 510874 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 511494 333978
rect 510874 316350 511494 333922
rect 510874 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 511494 316350
rect 510874 316226 511494 316294
rect 510874 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 511494 316226
rect 510874 316102 511494 316170
rect 510874 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 511494 316102
rect 510874 315978 511494 316046
rect 510874 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 511494 315978
rect 510874 298350 511494 315922
rect 510874 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 511494 298350
rect 510874 298226 511494 298294
rect 510874 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 511494 298226
rect 510874 298102 511494 298170
rect 510874 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 511494 298102
rect 510874 297978 511494 298046
rect 510874 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 511494 297978
rect 510874 280350 511494 297922
rect 510874 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 511494 280350
rect 510874 280226 511494 280294
rect 510874 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 511494 280226
rect 510874 280102 511494 280170
rect 510874 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 511494 280102
rect 510874 279978 511494 280046
rect 510874 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 511494 279978
rect 510874 262350 511494 279922
rect 510874 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 511494 262350
rect 510874 262226 511494 262294
rect 510874 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 511494 262226
rect 510874 262102 511494 262170
rect 510874 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 511494 262102
rect 510874 261978 511494 262046
rect 510874 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 511494 261978
rect 510874 244350 511494 261922
rect 510874 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 511494 244350
rect 510874 244226 511494 244294
rect 510874 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 511494 244226
rect 510874 244102 511494 244170
rect 510874 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 511494 244102
rect 510874 243978 511494 244046
rect 510874 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 511494 243978
rect 510874 226350 511494 243922
rect 510874 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 511494 226350
rect 510874 226226 511494 226294
rect 510874 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 511494 226226
rect 510874 226102 511494 226170
rect 510874 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 511494 226102
rect 510874 225978 511494 226046
rect 510874 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 511494 225978
rect 510874 208350 511494 225922
rect 510874 208294 510970 208350
rect 511026 208294 511094 208350
rect 511150 208294 511218 208350
rect 511274 208294 511342 208350
rect 511398 208294 511494 208350
rect 510874 208226 511494 208294
rect 510874 208170 510970 208226
rect 511026 208170 511094 208226
rect 511150 208170 511218 208226
rect 511274 208170 511342 208226
rect 511398 208170 511494 208226
rect 510874 208102 511494 208170
rect 510874 208046 510970 208102
rect 511026 208046 511094 208102
rect 511150 208046 511218 208102
rect 511274 208046 511342 208102
rect 511398 208046 511494 208102
rect 510874 207978 511494 208046
rect 510874 207922 510970 207978
rect 511026 207922 511094 207978
rect 511150 207922 511218 207978
rect 511274 207922 511342 207978
rect 511398 207922 511494 207978
rect 510874 190350 511494 207922
rect 510874 190294 510970 190350
rect 511026 190294 511094 190350
rect 511150 190294 511218 190350
rect 511274 190294 511342 190350
rect 511398 190294 511494 190350
rect 510874 190226 511494 190294
rect 510874 190170 510970 190226
rect 511026 190170 511094 190226
rect 511150 190170 511218 190226
rect 511274 190170 511342 190226
rect 511398 190170 511494 190226
rect 510874 190102 511494 190170
rect 510874 190046 510970 190102
rect 511026 190046 511094 190102
rect 511150 190046 511218 190102
rect 511274 190046 511342 190102
rect 511398 190046 511494 190102
rect 510874 189978 511494 190046
rect 510874 189922 510970 189978
rect 511026 189922 511094 189978
rect 511150 189922 511218 189978
rect 511274 189922 511342 189978
rect 511398 189922 511494 189978
rect 510874 172350 511494 189922
rect 510874 172294 510970 172350
rect 511026 172294 511094 172350
rect 511150 172294 511218 172350
rect 511274 172294 511342 172350
rect 511398 172294 511494 172350
rect 510874 172226 511494 172294
rect 510874 172170 510970 172226
rect 511026 172170 511094 172226
rect 511150 172170 511218 172226
rect 511274 172170 511342 172226
rect 511398 172170 511494 172226
rect 510874 172102 511494 172170
rect 510874 172046 510970 172102
rect 511026 172046 511094 172102
rect 511150 172046 511218 172102
rect 511274 172046 511342 172102
rect 511398 172046 511494 172102
rect 510874 171978 511494 172046
rect 510874 171922 510970 171978
rect 511026 171922 511094 171978
rect 511150 171922 511218 171978
rect 511274 171922 511342 171978
rect 511398 171922 511494 171978
rect 510874 154350 511494 171922
rect 510874 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 511494 154350
rect 510874 154226 511494 154294
rect 510874 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 511494 154226
rect 510874 154102 511494 154170
rect 510874 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 511494 154102
rect 510874 153978 511494 154046
rect 510874 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 511494 153978
rect 510874 136350 511494 153922
rect 510874 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 511494 136350
rect 510874 136226 511494 136294
rect 510874 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 511494 136226
rect 510874 136102 511494 136170
rect 510874 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 511494 136102
rect 510874 135978 511494 136046
rect 510874 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 511494 135978
rect 510874 118350 511494 135922
rect 510874 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 511494 118350
rect 510874 118226 511494 118294
rect 510874 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 511494 118226
rect 510874 118102 511494 118170
rect 510874 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 511494 118102
rect 510874 117978 511494 118046
rect 510874 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 511494 117978
rect 510874 100350 511494 117922
rect 510874 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 511494 100350
rect 510874 100226 511494 100294
rect 510874 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 511494 100226
rect 510874 100102 511494 100170
rect 510874 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 511494 100102
rect 510874 99978 511494 100046
rect 510874 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 511494 99978
rect 510874 82350 511494 99922
rect 510874 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 511494 82350
rect 510874 82226 511494 82294
rect 510874 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 511494 82226
rect 510874 82102 511494 82170
rect 510874 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 511494 82102
rect 510874 81978 511494 82046
rect 510874 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 511494 81978
rect 510874 64350 511494 81922
rect 510874 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 511494 64350
rect 510874 64226 511494 64294
rect 510874 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 511494 64226
rect 510874 64102 511494 64170
rect 510874 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 511494 64102
rect 510874 63978 511494 64046
rect 510874 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 511494 63978
rect 510874 46350 511494 63922
rect 510874 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 511494 46350
rect 510874 46226 511494 46294
rect 510874 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 511494 46226
rect 510874 46102 511494 46170
rect 510874 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 511494 46102
rect 510874 45978 511494 46046
rect 510874 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 511494 45978
rect 510874 28350 511494 45922
rect 510874 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 511494 28350
rect 510874 28226 511494 28294
rect 510874 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 511494 28226
rect 510874 28102 511494 28170
rect 510874 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 511494 28102
rect 510874 27978 511494 28046
rect 510874 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 511494 27978
rect 510874 10350 511494 27922
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 597212 525774 598268
rect 525154 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 525774 597212
rect 525154 597088 525774 597156
rect 525154 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 525774 597088
rect 525154 596964 525774 597032
rect 525154 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 525774 596964
rect 525154 596840 525774 596908
rect 525154 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 525774 596840
rect 525154 580350 525774 596784
rect 525154 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 525774 580350
rect 525154 580226 525774 580294
rect 525154 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 525774 580226
rect 525154 580102 525774 580170
rect 525154 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 525774 580102
rect 525154 579978 525774 580046
rect 525154 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 525774 579978
rect 525154 562350 525774 579922
rect 525154 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 525774 562350
rect 525154 562226 525774 562294
rect 525154 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 525774 562226
rect 525154 562102 525774 562170
rect 525154 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 525774 562102
rect 525154 561978 525774 562046
rect 525154 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 525774 561978
rect 525154 544350 525774 561922
rect 525154 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 525774 544350
rect 525154 544226 525774 544294
rect 525154 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 525774 544226
rect 525154 544102 525774 544170
rect 525154 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 525774 544102
rect 525154 543978 525774 544046
rect 525154 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 525774 543978
rect 525154 526350 525774 543922
rect 525154 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 525774 526350
rect 525154 526226 525774 526294
rect 525154 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 525774 526226
rect 525154 526102 525774 526170
rect 525154 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 525774 526102
rect 525154 525978 525774 526046
rect 525154 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 525774 525978
rect 525154 508350 525774 525922
rect 525154 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 525774 508350
rect 525154 508226 525774 508294
rect 525154 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 525774 508226
rect 525154 508102 525774 508170
rect 525154 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 525774 508102
rect 525154 507978 525774 508046
rect 525154 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 525774 507978
rect 525154 490350 525774 507922
rect 525154 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 525774 490350
rect 525154 490226 525774 490294
rect 525154 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 525774 490226
rect 525154 490102 525774 490170
rect 525154 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 525774 490102
rect 525154 489978 525774 490046
rect 525154 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 525774 489978
rect 525154 472350 525774 489922
rect 525154 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 525774 472350
rect 525154 472226 525774 472294
rect 525154 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 525774 472226
rect 525154 472102 525774 472170
rect 525154 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 525774 472102
rect 525154 471978 525774 472046
rect 525154 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 525774 471978
rect 525154 454350 525774 471922
rect 525154 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 525774 454350
rect 525154 454226 525774 454294
rect 525154 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 525774 454226
rect 525154 454102 525774 454170
rect 525154 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 525774 454102
rect 525154 453978 525774 454046
rect 525154 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 525774 453978
rect 525154 436350 525774 453922
rect 525154 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 525774 436350
rect 525154 436226 525774 436294
rect 525154 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 525774 436226
rect 525154 436102 525774 436170
rect 525154 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 525774 436102
rect 525154 435978 525774 436046
rect 525154 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 525774 435978
rect 525154 418350 525774 435922
rect 525154 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 525774 418350
rect 525154 418226 525774 418294
rect 525154 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 525774 418226
rect 525154 418102 525774 418170
rect 525154 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 525774 418102
rect 525154 417978 525774 418046
rect 525154 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 525774 417978
rect 525154 400350 525774 417922
rect 525154 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 525774 400350
rect 525154 400226 525774 400294
rect 525154 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 525774 400226
rect 525154 400102 525774 400170
rect 525154 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 525774 400102
rect 525154 399978 525774 400046
rect 525154 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 525774 399978
rect 525154 382350 525774 399922
rect 525154 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 525774 382350
rect 525154 382226 525774 382294
rect 525154 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 525774 382226
rect 525154 382102 525774 382170
rect 525154 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 525774 382102
rect 525154 381978 525774 382046
rect 525154 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 525774 381978
rect 525154 364350 525774 381922
rect 525154 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 525774 364350
rect 525154 364226 525774 364294
rect 525154 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 525774 364226
rect 525154 364102 525774 364170
rect 525154 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 525774 364102
rect 525154 363978 525774 364046
rect 525154 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 525774 363978
rect 525154 346350 525774 363922
rect 525154 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 525774 346350
rect 525154 346226 525774 346294
rect 525154 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 525774 346226
rect 525154 346102 525774 346170
rect 525154 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 525774 346102
rect 525154 345978 525774 346046
rect 525154 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 525774 345978
rect 525154 328350 525774 345922
rect 525154 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 525774 328350
rect 525154 328226 525774 328294
rect 525154 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 525774 328226
rect 525154 328102 525774 328170
rect 525154 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 525774 328102
rect 525154 327978 525774 328046
rect 525154 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 525774 327978
rect 525154 310350 525774 327922
rect 525154 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 525774 310350
rect 525154 310226 525774 310294
rect 525154 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 525774 310226
rect 525154 310102 525774 310170
rect 525154 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 525774 310102
rect 525154 309978 525774 310046
rect 525154 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 525774 309978
rect 525154 292350 525774 309922
rect 525154 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 525774 292350
rect 525154 292226 525774 292294
rect 525154 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 525774 292226
rect 525154 292102 525774 292170
rect 525154 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 525774 292102
rect 525154 291978 525774 292046
rect 525154 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 525774 291978
rect 525154 274350 525774 291922
rect 525154 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 525774 274350
rect 525154 274226 525774 274294
rect 525154 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 525774 274226
rect 525154 274102 525774 274170
rect 525154 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 525774 274102
rect 525154 273978 525774 274046
rect 525154 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 525774 273978
rect 525154 256350 525774 273922
rect 525154 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 525774 256350
rect 525154 256226 525774 256294
rect 525154 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 525774 256226
rect 525154 256102 525774 256170
rect 525154 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 525774 256102
rect 525154 255978 525774 256046
rect 525154 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 525774 255978
rect 525154 238350 525774 255922
rect 525154 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 525774 238350
rect 525154 238226 525774 238294
rect 525154 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 525774 238226
rect 525154 238102 525774 238170
rect 525154 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 525774 238102
rect 525154 237978 525774 238046
rect 525154 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 525774 237978
rect 525154 220350 525774 237922
rect 525154 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 525774 220350
rect 525154 220226 525774 220294
rect 525154 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 525774 220226
rect 525154 220102 525774 220170
rect 525154 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 525774 220102
rect 525154 219978 525774 220046
rect 525154 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 525774 219978
rect 525154 202350 525774 219922
rect 525154 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 525774 202350
rect 525154 202226 525774 202294
rect 525154 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 525774 202226
rect 525154 202102 525774 202170
rect 525154 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 525774 202102
rect 525154 201978 525774 202046
rect 525154 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 525774 201978
rect 525154 184350 525774 201922
rect 525154 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 525774 184350
rect 525154 184226 525774 184294
rect 525154 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 525774 184226
rect 525154 184102 525774 184170
rect 525154 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 525774 184102
rect 525154 183978 525774 184046
rect 525154 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 525774 183978
rect 525154 166350 525774 183922
rect 525154 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 525774 166350
rect 525154 166226 525774 166294
rect 525154 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 525774 166226
rect 525154 166102 525774 166170
rect 525154 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 525774 166102
rect 525154 165978 525774 166046
rect 525154 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 525774 165978
rect 525154 148350 525774 165922
rect 525154 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 525774 148350
rect 525154 148226 525774 148294
rect 525154 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 525774 148226
rect 525154 148102 525774 148170
rect 525154 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 525774 148102
rect 525154 147978 525774 148046
rect 525154 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 525774 147978
rect 525154 130350 525774 147922
rect 525154 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 525774 130350
rect 525154 130226 525774 130294
rect 525154 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 525774 130226
rect 525154 130102 525774 130170
rect 525154 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 525774 130102
rect 525154 129978 525774 130046
rect 525154 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 525774 129978
rect 525154 112350 525774 129922
rect 525154 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 525774 112350
rect 525154 112226 525774 112294
rect 525154 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 525774 112226
rect 525154 112102 525774 112170
rect 525154 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 525774 112102
rect 525154 111978 525774 112046
rect 525154 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 525774 111978
rect 525154 94350 525774 111922
rect 525154 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 525774 94350
rect 525154 94226 525774 94294
rect 525154 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 525774 94226
rect 525154 94102 525774 94170
rect 525154 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 525774 94102
rect 525154 93978 525774 94046
rect 525154 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 525774 93978
rect 525154 76350 525774 93922
rect 525154 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 525774 76350
rect 525154 76226 525774 76294
rect 525154 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 525774 76226
rect 525154 76102 525774 76170
rect 525154 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 525774 76102
rect 525154 75978 525774 76046
rect 525154 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 525774 75978
rect 525154 58350 525774 75922
rect 525154 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 525774 58350
rect 525154 58226 525774 58294
rect 525154 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 525774 58226
rect 525154 58102 525774 58170
rect 525154 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 525774 58102
rect 525154 57978 525774 58046
rect 525154 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 525774 57978
rect 525154 40350 525774 57922
rect 525154 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 525774 40350
rect 525154 40226 525774 40294
rect 525154 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 525774 40226
rect 525154 40102 525774 40170
rect 525154 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 525774 40102
rect 525154 39978 525774 40046
rect 525154 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 525774 39978
rect 525154 22350 525774 39922
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 514350 529494 531922
rect 528874 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 529494 514350
rect 528874 514226 529494 514294
rect 528874 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 529494 514226
rect 528874 514102 529494 514170
rect 528874 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 529494 514102
rect 528874 513978 529494 514046
rect 528874 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 529494 513978
rect 528874 496350 529494 513922
rect 528874 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 529494 496350
rect 528874 496226 529494 496294
rect 528874 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 529494 496226
rect 528874 496102 529494 496170
rect 528874 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 529494 496102
rect 528874 495978 529494 496046
rect 528874 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 529494 495978
rect 528874 478350 529494 495922
rect 528874 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 529494 478350
rect 528874 478226 529494 478294
rect 528874 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 529494 478226
rect 528874 478102 529494 478170
rect 528874 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 529494 478102
rect 528874 477978 529494 478046
rect 528874 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 529494 477978
rect 528874 460350 529494 477922
rect 528874 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 529494 460350
rect 528874 460226 529494 460294
rect 528874 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 529494 460226
rect 528874 460102 529494 460170
rect 528874 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 529494 460102
rect 528874 459978 529494 460046
rect 528874 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 529494 459978
rect 528874 442350 529494 459922
rect 528874 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 529494 442350
rect 528874 442226 529494 442294
rect 528874 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 529494 442226
rect 528874 442102 529494 442170
rect 528874 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 529494 442102
rect 528874 441978 529494 442046
rect 528874 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 529494 441978
rect 528874 424350 529494 441922
rect 528874 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 529494 424350
rect 528874 424226 529494 424294
rect 528874 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 529494 424226
rect 528874 424102 529494 424170
rect 528874 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 529494 424102
rect 528874 423978 529494 424046
rect 528874 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 529494 423978
rect 528874 406350 529494 423922
rect 528874 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 529494 406350
rect 528874 406226 529494 406294
rect 528874 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 529494 406226
rect 528874 406102 529494 406170
rect 528874 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 529494 406102
rect 528874 405978 529494 406046
rect 528874 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 529494 405978
rect 528874 388350 529494 405922
rect 528874 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 529494 388350
rect 528874 388226 529494 388294
rect 528874 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 529494 388226
rect 528874 388102 529494 388170
rect 528874 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 529494 388102
rect 528874 387978 529494 388046
rect 528874 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 529494 387978
rect 528874 370350 529494 387922
rect 528874 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 529494 370350
rect 528874 370226 529494 370294
rect 528874 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 529494 370226
rect 528874 370102 529494 370170
rect 528874 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 529494 370102
rect 528874 369978 529494 370046
rect 528874 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 529494 369978
rect 528874 352350 529494 369922
rect 528874 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 529494 352350
rect 528874 352226 529494 352294
rect 528874 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 529494 352226
rect 528874 352102 529494 352170
rect 528874 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 529494 352102
rect 528874 351978 529494 352046
rect 528874 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 529494 351978
rect 528874 334350 529494 351922
rect 528874 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 529494 334350
rect 528874 334226 529494 334294
rect 528874 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 529494 334226
rect 528874 334102 529494 334170
rect 528874 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 529494 334102
rect 528874 333978 529494 334046
rect 528874 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 529494 333978
rect 528874 316350 529494 333922
rect 528874 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 529494 316350
rect 528874 316226 529494 316294
rect 528874 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 529494 316226
rect 528874 316102 529494 316170
rect 528874 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 529494 316102
rect 528874 315978 529494 316046
rect 528874 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 529494 315978
rect 528874 298350 529494 315922
rect 528874 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 529494 298350
rect 528874 298226 529494 298294
rect 528874 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 529494 298226
rect 528874 298102 529494 298170
rect 528874 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 529494 298102
rect 528874 297978 529494 298046
rect 528874 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 529494 297978
rect 528874 280350 529494 297922
rect 528874 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 529494 280350
rect 528874 280226 529494 280294
rect 528874 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 529494 280226
rect 528874 280102 529494 280170
rect 528874 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 529494 280102
rect 528874 279978 529494 280046
rect 528874 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 529494 279978
rect 528874 262350 529494 279922
rect 528874 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 529494 262350
rect 528874 262226 529494 262294
rect 528874 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 529494 262226
rect 528874 262102 529494 262170
rect 528874 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 529494 262102
rect 528874 261978 529494 262046
rect 528874 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 529494 261978
rect 528874 244350 529494 261922
rect 528874 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 529494 244350
rect 528874 244226 529494 244294
rect 528874 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 529494 244226
rect 528874 244102 529494 244170
rect 528874 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 529494 244102
rect 528874 243978 529494 244046
rect 528874 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 529494 243978
rect 528874 226350 529494 243922
rect 528874 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 529494 226350
rect 528874 226226 529494 226294
rect 528874 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 529494 226226
rect 528874 226102 529494 226170
rect 528874 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 529494 226102
rect 528874 225978 529494 226046
rect 528874 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 529494 225978
rect 528874 208350 529494 225922
rect 528874 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 529494 208350
rect 528874 208226 529494 208294
rect 528874 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 529494 208226
rect 528874 208102 529494 208170
rect 528874 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 529494 208102
rect 528874 207978 529494 208046
rect 528874 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 529494 207978
rect 528874 190350 529494 207922
rect 528874 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 529494 190350
rect 528874 190226 529494 190294
rect 528874 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 529494 190226
rect 528874 190102 529494 190170
rect 528874 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 529494 190102
rect 528874 189978 529494 190046
rect 528874 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 529494 189978
rect 528874 172350 529494 189922
rect 528874 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 529494 172350
rect 528874 172226 529494 172294
rect 528874 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 529494 172226
rect 528874 172102 529494 172170
rect 528874 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 529494 172102
rect 528874 171978 529494 172046
rect 528874 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 529494 171978
rect 528874 154350 529494 171922
rect 528874 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 529494 154350
rect 528874 154226 529494 154294
rect 528874 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 529494 154226
rect 528874 154102 529494 154170
rect 528874 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 529494 154102
rect 528874 153978 529494 154046
rect 528874 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 529494 153978
rect 528874 136350 529494 153922
rect 528874 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 529494 136350
rect 528874 136226 529494 136294
rect 528874 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 529494 136226
rect 528874 136102 529494 136170
rect 528874 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 529494 136102
rect 528874 135978 529494 136046
rect 528874 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 529494 135978
rect 528874 118350 529494 135922
rect 528874 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 529494 118350
rect 528874 118226 529494 118294
rect 528874 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 529494 118226
rect 528874 118102 529494 118170
rect 528874 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 529494 118102
rect 528874 117978 529494 118046
rect 528874 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 529494 117978
rect 528874 100350 529494 117922
rect 528874 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 529494 100350
rect 528874 100226 529494 100294
rect 528874 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 529494 100226
rect 528874 100102 529494 100170
rect 528874 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 529494 100102
rect 528874 99978 529494 100046
rect 528874 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 529494 99978
rect 528874 82350 529494 99922
rect 528874 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 529494 82350
rect 528874 82226 529494 82294
rect 528874 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 529494 82226
rect 528874 82102 529494 82170
rect 528874 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 529494 82102
rect 528874 81978 529494 82046
rect 528874 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 529494 81978
rect 528874 64350 529494 81922
rect 528874 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 529494 64350
rect 528874 64226 529494 64294
rect 528874 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 529494 64226
rect 528874 64102 529494 64170
rect 528874 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 529494 64102
rect 528874 63978 529494 64046
rect 528874 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 529494 63978
rect 528874 46350 529494 63922
rect 528874 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 529494 46350
rect 528874 46226 529494 46294
rect 528874 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 529494 46226
rect 528874 46102 529494 46170
rect 528874 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 529494 46102
rect 528874 45978 529494 46046
rect 528874 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 529494 45978
rect 528874 28350 529494 45922
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 526350 543774 543922
rect 543154 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 543774 526350
rect 543154 526226 543774 526294
rect 543154 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 543774 526226
rect 543154 526102 543774 526170
rect 543154 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 543774 526102
rect 543154 525978 543774 526046
rect 543154 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 543774 525978
rect 543154 508350 543774 525922
rect 543154 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 543774 508350
rect 543154 508226 543774 508294
rect 543154 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 543774 508226
rect 543154 508102 543774 508170
rect 543154 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 543774 508102
rect 543154 507978 543774 508046
rect 543154 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 543774 507978
rect 543154 490350 543774 507922
rect 543154 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 543774 490350
rect 543154 490226 543774 490294
rect 543154 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 543774 490226
rect 543154 490102 543774 490170
rect 543154 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 543774 490102
rect 543154 489978 543774 490046
rect 543154 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 543774 489978
rect 543154 472350 543774 489922
rect 543154 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 543774 472350
rect 543154 472226 543774 472294
rect 543154 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 543774 472226
rect 543154 472102 543774 472170
rect 543154 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 543774 472102
rect 543154 471978 543774 472046
rect 543154 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 543774 471978
rect 543154 454350 543774 471922
rect 543154 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 543774 454350
rect 543154 454226 543774 454294
rect 543154 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 543774 454226
rect 543154 454102 543774 454170
rect 543154 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 543774 454102
rect 543154 453978 543774 454046
rect 543154 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 543774 453978
rect 543154 436350 543774 453922
rect 543154 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 543774 436350
rect 543154 436226 543774 436294
rect 543154 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 543774 436226
rect 543154 436102 543774 436170
rect 543154 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 543774 436102
rect 543154 435978 543774 436046
rect 543154 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 543774 435978
rect 543154 418350 543774 435922
rect 543154 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 543774 418350
rect 543154 418226 543774 418294
rect 543154 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 543774 418226
rect 543154 418102 543774 418170
rect 543154 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 543774 418102
rect 543154 417978 543774 418046
rect 543154 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 543774 417978
rect 543154 400350 543774 417922
rect 543154 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 543774 400350
rect 543154 400226 543774 400294
rect 543154 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 543774 400226
rect 543154 400102 543774 400170
rect 543154 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 543774 400102
rect 543154 399978 543774 400046
rect 543154 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 543774 399978
rect 543154 382350 543774 399922
rect 543154 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 543774 382350
rect 543154 382226 543774 382294
rect 543154 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 543774 382226
rect 543154 382102 543774 382170
rect 543154 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 543774 382102
rect 543154 381978 543774 382046
rect 543154 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 543774 381978
rect 543154 364350 543774 381922
rect 543154 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 543774 364350
rect 543154 364226 543774 364294
rect 543154 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 543774 364226
rect 543154 364102 543774 364170
rect 543154 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 543774 364102
rect 543154 363978 543774 364046
rect 543154 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 543774 363978
rect 543154 346350 543774 363922
rect 543154 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 543774 346350
rect 543154 346226 543774 346294
rect 543154 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 543774 346226
rect 543154 346102 543774 346170
rect 543154 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 543774 346102
rect 543154 345978 543774 346046
rect 543154 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 543774 345978
rect 543154 328350 543774 345922
rect 543154 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 543774 328350
rect 543154 328226 543774 328294
rect 543154 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 543774 328226
rect 543154 328102 543774 328170
rect 543154 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 543774 328102
rect 543154 327978 543774 328046
rect 543154 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 543774 327978
rect 543154 310350 543774 327922
rect 543154 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 543774 310350
rect 543154 310226 543774 310294
rect 543154 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 543774 310226
rect 543154 310102 543774 310170
rect 543154 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 543774 310102
rect 543154 309978 543774 310046
rect 543154 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 543774 309978
rect 543154 292350 543774 309922
rect 543154 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 543774 292350
rect 543154 292226 543774 292294
rect 543154 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 543774 292226
rect 543154 292102 543774 292170
rect 543154 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 543774 292102
rect 543154 291978 543774 292046
rect 543154 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 543774 291978
rect 543154 274350 543774 291922
rect 543154 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 543774 274350
rect 543154 274226 543774 274294
rect 543154 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 543774 274226
rect 543154 274102 543774 274170
rect 543154 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 543774 274102
rect 543154 273978 543774 274046
rect 543154 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 543774 273978
rect 543154 256350 543774 273922
rect 543154 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 543774 256350
rect 543154 256226 543774 256294
rect 543154 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 543774 256226
rect 543154 256102 543774 256170
rect 543154 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 543774 256102
rect 543154 255978 543774 256046
rect 543154 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 543774 255978
rect 543154 238350 543774 255922
rect 543154 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 543774 238350
rect 543154 238226 543774 238294
rect 543154 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 543774 238226
rect 543154 238102 543774 238170
rect 543154 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 543774 238102
rect 543154 237978 543774 238046
rect 543154 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 543774 237978
rect 543154 220350 543774 237922
rect 543154 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 543774 220350
rect 543154 220226 543774 220294
rect 543154 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 543774 220226
rect 543154 220102 543774 220170
rect 543154 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 543774 220102
rect 543154 219978 543774 220046
rect 543154 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 543774 219978
rect 543154 202350 543774 219922
rect 543154 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 543774 202350
rect 543154 202226 543774 202294
rect 543154 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 543774 202226
rect 543154 202102 543774 202170
rect 543154 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 543774 202102
rect 543154 201978 543774 202046
rect 543154 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 543774 201978
rect 543154 184350 543774 201922
rect 543154 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 543774 184350
rect 543154 184226 543774 184294
rect 543154 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 543774 184226
rect 543154 184102 543774 184170
rect 543154 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 543774 184102
rect 543154 183978 543774 184046
rect 543154 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 543774 183978
rect 543154 166350 543774 183922
rect 543154 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 543774 166350
rect 543154 166226 543774 166294
rect 543154 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 543774 166226
rect 543154 166102 543774 166170
rect 543154 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 543774 166102
rect 543154 165978 543774 166046
rect 543154 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 543774 165978
rect 543154 148350 543774 165922
rect 543154 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 543774 148350
rect 543154 148226 543774 148294
rect 543154 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 543774 148226
rect 543154 148102 543774 148170
rect 543154 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 543774 148102
rect 543154 147978 543774 148046
rect 543154 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 543774 147978
rect 543154 130350 543774 147922
rect 543154 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 543774 130350
rect 543154 130226 543774 130294
rect 543154 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 543774 130226
rect 543154 130102 543774 130170
rect 543154 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 543774 130102
rect 543154 129978 543774 130046
rect 543154 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 543774 129978
rect 543154 112350 543774 129922
rect 543154 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 543774 112350
rect 543154 112226 543774 112294
rect 543154 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 543774 112226
rect 543154 112102 543774 112170
rect 543154 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 543774 112102
rect 543154 111978 543774 112046
rect 543154 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 543774 111978
rect 543154 94350 543774 111922
rect 543154 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 543774 94350
rect 543154 94226 543774 94294
rect 543154 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 543774 94226
rect 543154 94102 543774 94170
rect 543154 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 543774 94102
rect 543154 93978 543774 94046
rect 543154 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 543774 93978
rect 543154 76350 543774 93922
rect 543154 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 543774 76350
rect 543154 76226 543774 76294
rect 543154 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 543774 76226
rect 543154 76102 543774 76170
rect 543154 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 543774 76102
rect 543154 75978 543774 76046
rect 543154 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 543774 75978
rect 543154 58350 543774 75922
rect 543154 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 543774 58350
rect 543154 58226 543774 58294
rect 543154 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 543774 58226
rect 543154 58102 543774 58170
rect 543154 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 543774 58102
rect 543154 57978 543774 58046
rect 543154 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 543774 57978
rect 543154 40350 543774 57922
rect 543154 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 543774 40350
rect 543154 40226 543774 40294
rect 543154 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 543774 40226
rect 543154 40102 543774 40170
rect 543154 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 543774 40102
rect 543154 39978 543774 40046
rect 543154 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 543774 39978
rect 543154 22350 543774 39922
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 514350 547494 531922
rect 546874 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 547494 514350
rect 546874 514226 547494 514294
rect 546874 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 547494 514226
rect 546874 514102 547494 514170
rect 546874 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 547494 514102
rect 546874 513978 547494 514046
rect 546874 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 547494 513978
rect 546874 496350 547494 513922
rect 546874 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 547494 496350
rect 546874 496226 547494 496294
rect 546874 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 547494 496226
rect 546874 496102 547494 496170
rect 546874 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 547494 496102
rect 546874 495978 547494 496046
rect 546874 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 547494 495978
rect 546874 478350 547494 495922
rect 546874 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 547494 478350
rect 546874 478226 547494 478294
rect 546874 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 547494 478226
rect 546874 478102 547494 478170
rect 546874 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 547494 478102
rect 546874 477978 547494 478046
rect 546874 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 547494 477978
rect 546874 460350 547494 477922
rect 546874 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 547494 460350
rect 546874 460226 547494 460294
rect 546874 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 547494 460226
rect 546874 460102 547494 460170
rect 546874 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 547494 460102
rect 546874 459978 547494 460046
rect 546874 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 547494 459978
rect 546874 442350 547494 459922
rect 546874 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 547494 442350
rect 546874 442226 547494 442294
rect 546874 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 547494 442226
rect 546874 442102 547494 442170
rect 546874 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 547494 442102
rect 546874 441978 547494 442046
rect 546874 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 547494 441978
rect 546874 424350 547494 441922
rect 546874 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 547494 424350
rect 546874 424226 547494 424294
rect 546874 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 547494 424226
rect 546874 424102 547494 424170
rect 546874 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 547494 424102
rect 546874 423978 547494 424046
rect 546874 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 547494 423978
rect 546874 406350 547494 423922
rect 546874 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 547494 406350
rect 546874 406226 547494 406294
rect 546874 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 547494 406226
rect 546874 406102 547494 406170
rect 546874 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 547494 406102
rect 546874 405978 547494 406046
rect 546874 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 547494 405978
rect 546874 388350 547494 405922
rect 546874 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 547494 388350
rect 546874 388226 547494 388294
rect 546874 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 547494 388226
rect 546874 388102 547494 388170
rect 546874 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 547494 388102
rect 546874 387978 547494 388046
rect 546874 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 547494 387978
rect 546874 370350 547494 387922
rect 546874 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 547494 370350
rect 546874 370226 547494 370294
rect 546874 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 547494 370226
rect 546874 370102 547494 370170
rect 546874 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 547494 370102
rect 546874 369978 547494 370046
rect 546874 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 547494 369978
rect 546874 352350 547494 369922
rect 546874 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 547494 352350
rect 546874 352226 547494 352294
rect 546874 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 547494 352226
rect 546874 352102 547494 352170
rect 546874 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 547494 352102
rect 546874 351978 547494 352046
rect 546874 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 547494 351978
rect 546874 334350 547494 351922
rect 546874 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 547494 334350
rect 546874 334226 547494 334294
rect 546874 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 547494 334226
rect 546874 334102 547494 334170
rect 546874 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 547494 334102
rect 546874 333978 547494 334046
rect 546874 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 547494 333978
rect 546874 316350 547494 333922
rect 546874 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 547494 316350
rect 546874 316226 547494 316294
rect 546874 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 547494 316226
rect 546874 316102 547494 316170
rect 546874 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 547494 316102
rect 546874 315978 547494 316046
rect 546874 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 547494 315978
rect 546874 298350 547494 315922
rect 546874 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 547494 298350
rect 546874 298226 547494 298294
rect 546874 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 547494 298226
rect 546874 298102 547494 298170
rect 546874 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 547494 298102
rect 546874 297978 547494 298046
rect 546874 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 547494 297978
rect 546874 280350 547494 297922
rect 546874 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 547494 280350
rect 546874 280226 547494 280294
rect 546874 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 547494 280226
rect 546874 280102 547494 280170
rect 546874 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 547494 280102
rect 546874 279978 547494 280046
rect 546874 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 547494 279978
rect 546874 262350 547494 279922
rect 546874 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 547494 262350
rect 546874 262226 547494 262294
rect 546874 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 547494 262226
rect 546874 262102 547494 262170
rect 546874 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 547494 262102
rect 546874 261978 547494 262046
rect 546874 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 547494 261978
rect 546874 244350 547494 261922
rect 546874 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 547494 244350
rect 546874 244226 547494 244294
rect 546874 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 547494 244226
rect 546874 244102 547494 244170
rect 546874 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 547494 244102
rect 546874 243978 547494 244046
rect 546874 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 547494 243978
rect 546874 226350 547494 243922
rect 546874 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 547494 226350
rect 546874 226226 547494 226294
rect 546874 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 547494 226226
rect 546874 226102 547494 226170
rect 546874 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 547494 226102
rect 546874 225978 547494 226046
rect 546874 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 547494 225978
rect 546874 208350 547494 225922
rect 546874 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 547494 208350
rect 546874 208226 547494 208294
rect 546874 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 547494 208226
rect 546874 208102 547494 208170
rect 546874 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 547494 208102
rect 546874 207978 547494 208046
rect 546874 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 547494 207978
rect 546874 190350 547494 207922
rect 546874 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 547494 190350
rect 546874 190226 547494 190294
rect 546874 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 547494 190226
rect 546874 190102 547494 190170
rect 546874 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 547494 190102
rect 546874 189978 547494 190046
rect 546874 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 547494 189978
rect 546874 172350 547494 189922
rect 546874 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 547494 172350
rect 546874 172226 547494 172294
rect 546874 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 547494 172226
rect 546874 172102 547494 172170
rect 546874 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 547494 172102
rect 546874 171978 547494 172046
rect 546874 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 547494 171978
rect 546874 154350 547494 171922
rect 546874 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 547494 154350
rect 546874 154226 547494 154294
rect 546874 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 547494 154226
rect 546874 154102 547494 154170
rect 546874 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 547494 154102
rect 546874 153978 547494 154046
rect 546874 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 547494 153978
rect 546874 136350 547494 153922
rect 546874 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 547494 136350
rect 546874 136226 547494 136294
rect 546874 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 547494 136226
rect 546874 136102 547494 136170
rect 546874 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 547494 136102
rect 546874 135978 547494 136046
rect 546874 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 547494 135978
rect 546874 118350 547494 135922
rect 546874 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 547494 118350
rect 546874 118226 547494 118294
rect 546874 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 547494 118226
rect 546874 118102 547494 118170
rect 546874 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 547494 118102
rect 546874 117978 547494 118046
rect 546874 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 547494 117978
rect 546874 100350 547494 117922
rect 546874 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 547494 100350
rect 546874 100226 547494 100294
rect 546874 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 547494 100226
rect 546874 100102 547494 100170
rect 546874 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 547494 100102
rect 546874 99978 547494 100046
rect 546874 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 547494 99978
rect 546874 82350 547494 99922
rect 546874 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 547494 82350
rect 546874 82226 547494 82294
rect 546874 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 547494 82226
rect 546874 82102 547494 82170
rect 546874 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 547494 82102
rect 546874 81978 547494 82046
rect 546874 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 547494 81978
rect 546874 64350 547494 81922
rect 546874 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 547494 64350
rect 546874 64226 547494 64294
rect 546874 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 547494 64226
rect 546874 64102 547494 64170
rect 546874 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 547494 64102
rect 546874 63978 547494 64046
rect 546874 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 547494 63978
rect 546874 46350 547494 63922
rect 546874 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 547494 46350
rect 546874 46226 547494 46294
rect 546874 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 547494 46226
rect 546874 46102 547494 46170
rect 546874 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 547494 46102
rect 546874 45978 547494 46046
rect 546874 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 547494 45978
rect 546874 28350 547494 45922
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 561154 526350 561774 543922
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 561154 490350 561774 507922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 561154 472350 561774 489922
rect 561154 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 561774 472350
rect 561154 472226 561774 472294
rect 561154 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 561774 472226
rect 561154 472102 561774 472170
rect 561154 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 561774 472102
rect 561154 471978 561774 472046
rect 561154 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 561774 471978
rect 561154 454350 561774 471922
rect 561154 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 561774 454350
rect 561154 454226 561774 454294
rect 561154 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 561774 454226
rect 561154 454102 561774 454170
rect 561154 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 561774 454102
rect 561154 453978 561774 454046
rect 561154 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 561774 453978
rect 561154 436350 561774 453922
rect 561154 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 561774 436350
rect 561154 436226 561774 436294
rect 561154 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 561774 436226
rect 561154 436102 561774 436170
rect 561154 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 561774 436102
rect 561154 435978 561774 436046
rect 561154 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 561774 435978
rect 561154 418350 561774 435922
rect 561154 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 561774 418350
rect 561154 418226 561774 418294
rect 561154 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 561774 418226
rect 561154 418102 561774 418170
rect 561154 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 561774 418102
rect 561154 417978 561774 418046
rect 561154 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 561774 417978
rect 561154 400350 561774 417922
rect 561154 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 561774 400350
rect 561154 400226 561774 400294
rect 561154 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 561774 400226
rect 561154 400102 561774 400170
rect 561154 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 561774 400102
rect 561154 399978 561774 400046
rect 561154 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 561774 399978
rect 561154 382350 561774 399922
rect 561154 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 561774 382350
rect 561154 382226 561774 382294
rect 561154 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 561774 382226
rect 561154 382102 561774 382170
rect 561154 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 561774 382102
rect 561154 381978 561774 382046
rect 561154 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 561774 381978
rect 561154 364350 561774 381922
rect 561154 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 561774 364350
rect 561154 364226 561774 364294
rect 561154 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 561774 364226
rect 561154 364102 561774 364170
rect 561154 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 561774 364102
rect 561154 363978 561774 364046
rect 561154 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 561774 363978
rect 561154 346350 561774 363922
rect 561154 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 561774 346350
rect 561154 346226 561774 346294
rect 561154 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 561774 346226
rect 561154 346102 561774 346170
rect 561154 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 561774 346102
rect 561154 345978 561774 346046
rect 561154 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 561774 345978
rect 561154 328350 561774 345922
rect 561154 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 561774 328350
rect 561154 328226 561774 328294
rect 561154 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 561774 328226
rect 561154 328102 561774 328170
rect 561154 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 561774 328102
rect 561154 327978 561774 328046
rect 561154 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 561774 327978
rect 561154 310350 561774 327922
rect 561154 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 561774 310350
rect 561154 310226 561774 310294
rect 561154 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 561774 310226
rect 561154 310102 561774 310170
rect 561154 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 561774 310102
rect 561154 309978 561774 310046
rect 561154 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 561774 309978
rect 561154 292350 561774 309922
rect 561154 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 561774 292350
rect 561154 292226 561774 292294
rect 561154 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 561774 292226
rect 561154 292102 561774 292170
rect 561154 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 561774 292102
rect 561154 291978 561774 292046
rect 561154 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 561774 291978
rect 561154 274350 561774 291922
rect 561154 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 561774 274350
rect 561154 274226 561774 274294
rect 561154 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 561774 274226
rect 561154 274102 561774 274170
rect 561154 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 561774 274102
rect 561154 273978 561774 274046
rect 561154 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 561774 273978
rect 561154 256350 561774 273922
rect 561154 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 561774 256350
rect 561154 256226 561774 256294
rect 561154 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 561774 256226
rect 561154 256102 561774 256170
rect 561154 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 561774 256102
rect 561154 255978 561774 256046
rect 561154 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 561774 255978
rect 561154 238350 561774 255922
rect 561154 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 561774 238350
rect 561154 238226 561774 238294
rect 561154 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 561774 238226
rect 561154 238102 561774 238170
rect 561154 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 561774 238102
rect 561154 237978 561774 238046
rect 561154 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 561774 237978
rect 561154 220350 561774 237922
rect 561154 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 561774 220350
rect 561154 220226 561774 220294
rect 561154 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 561774 220226
rect 561154 220102 561774 220170
rect 561154 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 561774 220102
rect 561154 219978 561774 220046
rect 561154 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 561774 219978
rect 561154 202350 561774 219922
rect 561154 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 561774 202350
rect 561154 202226 561774 202294
rect 561154 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 561774 202226
rect 561154 202102 561774 202170
rect 561154 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 561774 202102
rect 561154 201978 561774 202046
rect 561154 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 561774 201978
rect 561154 184350 561774 201922
rect 561154 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 561774 184350
rect 561154 184226 561774 184294
rect 561154 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 561774 184226
rect 561154 184102 561774 184170
rect 561154 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 561774 184102
rect 561154 183978 561774 184046
rect 561154 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 561774 183978
rect 561154 166350 561774 183922
rect 561154 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 561774 166350
rect 561154 166226 561774 166294
rect 561154 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 561774 166226
rect 561154 166102 561774 166170
rect 561154 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 561774 166102
rect 561154 165978 561774 166046
rect 561154 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 561774 165978
rect 561154 148350 561774 165922
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 561154 130350 561774 147922
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 561154 40350 561774 57922
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 561154 22350 561774 39922
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 4350 561774 21922
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 561154 -160 561774 3922
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 496350 565494 513922
rect 564874 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 565494 496350
rect 564874 496226 565494 496294
rect 564874 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 565494 496226
rect 564874 496102 565494 496170
rect 564874 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 565494 496102
rect 564874 495978 565494 496046
rect 564874 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 565494 495978
rect 564874 478350 565494 495922
rect 564874 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 565494 478350
rect 564874 478226 565494 478294
rect 564874 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 565494 478226
rect 564874 478102 565494 478170
rect 564874 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 565494 478102
rect 564874 477978 565494 478046
rect 564874 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 565494 477978
rect 564874 460350 565494 477922
rect 564874 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 565494 460350
rect 564874 460226 565494 460294
rect 564874 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 565494 460226
rect 564874 460102 565494 460170
rect 564874 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 565494 460102
rect 564874 459978 565494 460046
rect 564874 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 565494 459978
rect 564874 442350 565494 459922
rect 564874 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 565494 442350
rect 564874 442226 565494 442294
rect 564874 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 565494 442226
rect 564874 442102 565494 442170
rect 564874 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 565494 442102
rect 564874 441978 565494 442046
rect 564874 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 565494 441978
rect 564874 424350 565494 441922
rect 564874 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 565494 424350
rect 564874 424226 565494 424294
rect 564874 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 565494 424226
rect 564874 424102 565494 424170
rect 564874 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 565494 424102
rect 564874 423978 565494 424046
rect 564874 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 565494 423978
rect 564874 406350 565494 423922
rect 564874 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 565494 406350
rect 564874 406226 565494 406294
rect 564874 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 565494 406226
rect 564874 406102 565494 406170
rect 564874 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 565494 406102
rect 564874 405978 565494 406046
rect 564874 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 565494 405978
rect 564874 388350 565494 405922
rect 564874 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 565494 388350
rect 564874 388226 565494 388294
rect 564874 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 565494 388226
rect 564874 388102 565494 388170
rect 564874 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 565494 388102
rect 564874 387978 565494 388046
rect 564874 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 565494 387978
rect 564874 370350 565494 387922
rect 564874 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 565494 370350
rect 564874 370226 565494 370294
rect 564874 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 565494 370226
rect 564874 370102 565494 370170
rect 564874 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 565494 370102
rect 564874 369978 565494 370046
rect 564874 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 565494 369978
rect 564874 352350 565494 369922
rect 564874 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 565494 352350
rect 564874 352226 565494 352294
rect 564874 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 565494 352226
rect 564874 352102 565494 352170
rect 564874 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 565494 352102
rect 564874 351978 565494 352046
rect 564874 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 565494 351978
rect 564874 334350 565494 351922
rect 564874 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 565494 334350
rect 564874 334226 565494 334294
rect 564874 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 565494 334226
rect 564874 334102 565494 334170
rect 564874 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 565494 334102
rect 564874 333978 565494 334046
rect 564874 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 565494 333978
rect 564874 316350 565494 333922
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298350 565494 315922
rect 564874 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 565494 298350
rect 564874 298226 565494 298294
rect 564874 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 565494 298226
rect 564874 298102 565494 298170
rect 564874 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 565494 298102
rect 564874 297978 565494 298046
rect 564874 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 565494 297978
rect 564874 280350 565494 297922
rect 564874 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 565494 280350
rect 564874 280226 565494 280294
rect 564874 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 565494 280226
rect 564874 280102 565494 280170
rect 564874 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 565494 280102
rect 564874 279978 565494 280046
rect 564874 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 565494 279978
rect 564874 262350 565494 279922
rect 564874 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 565494 262350
rect 564874 262226 565494 262294
rect 564874 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 565494 262226
rect 564874 262102 565494 262170
rect 564874 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 565494 262102
rect 564874 261978 565494 262046
rect 564874 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 565494 261978
rect 564874 244350 565494 261922
rect 564874 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 565494 244350
rect 564874 244226 565494 244294
rect 564874 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 565494 244226
rect 564874 244102 565494 244170
rect 564874 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 565494 244102
rect 564874 243978 565494 244046
rect 564874 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 565494 243978
rect 564874 226350 565494 243922
rect 564874 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 565494 226350
rect 564874 226226 565494 226294
rect 564874 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 565494 226226
rect 564874 226102 565494 226170
rect 564874 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 565494 226102
rect 564874 225978 565494 226046
rect 564874 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 565494 225978
rect 564874 208350 565494 225922
rect 564874 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 565494 208350
rect 564874 208226 565494 208294
rect 564874 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 565494 208226
rect 564874 208102 565494 208170
rect 564874 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 565494 208102
rect 564874 207978 565494 208046
rect 564874 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 565494 207978
rect 564874 190350 565494 207922
rect 564874 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 565494 190350
rect 564874 190226 565494 190294
rect 564874 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 565494 190226
rect 564874 190102 565494 190170
rect 564874 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 565494 190102
rect 564874 189978 565494 190046
rect 564874 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 565494 189978
rect 564874 172350 565494 189922
rect 564874 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 565494 172350
rect 564874 172226 565494 172294
rect 564874 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 565494 172226
rect 564874 172102 565494 172170
rect 564874 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 565494 172102
rect 564874 171978 565494 172046
rect 564874 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 565494 171978
rect 564874 154350 565494 171922
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 564874 28350 565494 45922
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 10350 565494 27922
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 564874 -1120 565494 9922
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 579154 490350 579774 507922
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 472350 579774 489922
rect 579154 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 579774 472350
rect 579154 472226 579774 472294
rect 579154 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 579774 472226
rect 579154 472102 579774 472170
rect 579154 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 579774 472102
rect 579154 471978 579774 472046
rect 579154 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 579774 471978
rect 579154 454350 579774 471922
rect 579154 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 579774 454350
rect 579154 454226 579774 454294
rect 579154 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 579774 454226
rect 579154 454102 579774 454170
rect 579154 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 579774 454102
rect 579154 453978 579774 454046
rect 579154 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 579774 453978
rect 579154 436350 579774 453922
rect 579154 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 579774 436350
rect 579154 436226 579774 436294
rect 579154 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 579774 436226
rect 579154 436102 579774 436170
rect 579154 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 579774 436102
rect 579154 435978 579774 436046
rect 579154 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 579774 435978
rect 579154 418350 579774 435922
rect 579154 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 579774 418350
rect 579154 418226 579774 418294
rect 579154 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 579774 418226
rect 579154 418102 579774 418170
rect 579154 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 579774 418102
rect 579154 417978 579774 418046
rect 579154 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 579774 417978
rect 579154 400350 579774 417922
rect 579154 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 579774 400350
rect 579154 400226 579774 400294
rect 579154 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 579774 400226
rect 579154 400102 579774 400170
rect 579154 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 579774 400102
rect 579154 399978 579774 400046
rect 579154 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 579774 399978
rect 579154 382350 579774 399922
rect 579154 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 579774 382350
rect 579154 382226 579774 382294
rect 579154 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 579774 382226
rect 579154 382102 579774 382170
rect 579154 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 579774 382102
rect 579154 381978 579774 382046
rect 579154 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 579774 381978
rect 579154 364350 579774 381922
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58350 579774 75922
rect 579154 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 579774 58350
rect 579154 58226 579774 58294
rect 579154 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 579774 58226
rect 579154 58102 579774 58170
rect 579154 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 579774 58102
rect 579154 57978 579774 58046
rect 579154 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 579774 57978
rect 579154 40350 579774 57922
rect 579154 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 579774 40350
rect 579154 40226 579774 40294
rect 579154 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 579774 40226
rect 579154 40102 579774 40170
rect 579154 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 579774 40102
rect 579154 39978 579774 40046
rect 579154 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 579774 39978
rect 579154 22350 579774 39922
rect 579154 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 579774 22350
rect 579154 22226 579774 22294
rect 579154 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 579774 22226
rect 579154 22102 579774 22170
rect 579154 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 579774 22102
rect 579154 21978 579774 22046
rect 579154 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 579774 21978
rect 579154 4350 579774 21922
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 582874 496350 583494 513922
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 582874 478350 583494 495922
rect 582874 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 583494 478350
rect 582874 478226 583494 478294
rect 582874 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 583494 478226
rect 582874 478102 583494 478170
rect 582874 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 583494 478102
rect 582874 477978 583494 478046
rect 582874 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 583494 477978
rect 582874 460350 583494 477922
rect 582874 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 583494 460350
rect 582874 460226 583494 460294
rect 582874 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 583494 460226
rect 582874 460102 583494 460170
rect 582874 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 583494 460102
rect 582874 459978 583494 460046
rect 582874 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 583494 459978
rect 582874 442350 583494 459922
rect 582874 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 583494 442350
rect 582874 442226 583494 442294
rect 582874 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 583494 442226
rect 582874 442102 583494 442170
rect 582874 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 583494 442102
rect 582874 441978 583494 442046
rect 582874 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 583494 441978
rect 582874 424350 583494 441922
rect 582874 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 583494 424350
rect 582874 424226 583494 424294
rect 582874 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 583494 424226
rect 582874 424102 583494 424170
rect 582874 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 583494 424102
rect 582874 423978 583494 424046
rect 582874 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 583494 423978
rect 582874 406350 583494 423922
rect 582874 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 583494 406350
rect 582874 406226 583494 406294
rect 582874 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 583494 406226
rect 582874 406102 583494 406170
rect 582874 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 583494 406102
rect 582874 405978 583494 406046
rect 582874 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 583494 405978
rect 582874 388350 583494 405922
rect 582874 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 583494 388350
rect 582874 388226 583494 388294
rect 582874 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 583494 388226
rect 582874 388102 583494 388170
rect 582874 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 583494 388102
rect 582874 387978 583494 388046
rect 582874 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 583494 387978
rect 582874 370350 583494 387922
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 582874 -1120 583494 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 21250 508294 21306 508350
rect 21374 508294 21430 508350
rect 21498 508294 21554 508350
rect 21622 508294 21678 508350
rect 21250 508170 21306 508226
rect 21374 508170 21430 508226
rect 21498 508170 21554 508226
rect 21622 508170 21678 508226
rect 21250 508046 21306 508102
rect 21374 508046 21430 508102
rect 21498 508046 21554 508102
rect 21622 508046 21678 508102
rect 21250 507922 21306 507978
rect 21374 507922 21430 507978
rect 21498 507922 21554 507978
rect 21622 507922 21678 507978
rect 21250 490294 21306 490350
rect 21374 490294 21430 490350
rect 21498 490294 21554 490350
rect 21622 490294 21678 490350
rect 21250 490170 21306 490226
rect 21374 490170 21430 490226
rect 21498 490170 21554 490226
rect 21622 490170 21678 490226
rect 21250 490046 21306 490102
rect 21374 490046 21430 490102
rect 21498 490046 21554 490102
rect 21622 490046 21678 490102
rect 21250 489922 21306 489978
rect 21374 489922 21430 489978
rect 21498 489922 21554 489978
rect 21622 489922 21678 489978
rect 21250 472294 21306 472350
rect 21374 472294 21430 472350
rect 21498 472294 21554 472350
rect 21622 472294 21678 472350
rect 21250 472170 21306 472226
rect 21374 472170 21430 472226
rect 21498 472170 21554 472226
rect 21622 472170 21678 472226
rect 21250 472046 21306 472102
rect 21374 472046 21430 472102
rect 21498 472046 21554 472102
rect 21622 472046 21678 472102
rect 21250 471922 21306 471978
rect 21374 471922 21430 471978
rect 21498 471922 21554 471978
rect 21622 471922 21678 471978
rect 21250 454294 21306 454350
rect 21374 454294 21430 454350
rect 21498 454294 21554 454350
rect 21622 454294 21678 454350
rect 21250 454170 21306 454226
rect 21374 454170 21430 454226
rect 21498 454170 21554 454226
rect 21622 454170 21678 454226
rect 21250 454046 21306 454102
rect 21374 454046 21430 454102
rect 21498 454046 21554 454102
rect 21622 454046 21678 454102
rect 21250 453922 21306 453978
rect 21374 453922 21430 453978
rect 21498 453922 21554 453978
rect 21622 453922 21678 453978
rect 21250 436294 21306 436350
rect 21374 436294 21430 436350
rect 21498 436294 21554 436350
rect 21622 436294 21678 436350
rect 21250 436170 21306 436226
rect 21374 436170 21430 436226
rect 21498 436170 21554 436226
rect 21622 436170 21678 436226
rect 21250 436046 21306 436102
rect 21374 436046 21430 436102
rect 21498 436046 21554 436102
rect 21622 436046 21678 436102
rect 21250 435922 21306 435978
rect 21374 435922 21430 435978
rect 21498 435922 21554 435978
rect 21622 435922 21678 435978
rect 21250 418294 21306 418350
rect 21374 418294 21430 418350
rect 21498 418294 21554 418350
rect 21622 418294 21678 418350
rect 21250 418170 21306 418226
rect 21374 418170 21430 418226
rect 21498 418170 21554 418226
rect 21622 418170 21678 418226
rect 21250 418046 21306 418102
rect 21374 418046 21430 418102
rect 21498 418046 21554 418102
rect 21622 418046 21678 418102
rect 21250 417922 21306 417978
rect 21374 417922 21430 417978
rect 21498 417922 21554 417978
rect 21622 417922 21678 417978
rect 21250 400294 21306 400350
rect 21374 400294 21430 400350
rect 21498 400294 21554 400350
rect 21622 400294 21678 400350
rect 21250 400170 21306 400226
rect 21374 400170 21430 400226
rect 21498 400170 21554 400226
rect 21622 400170 21678 400226
rect 21250 400046 21306 400102
rect 21374 400046 21430 400102
rect 21498 400046 21554 400102
rect 21622 400046 21678 400102
rect 21250 399922 21306 399978
rect 21374 399922 21430 399978
rect 21498 399922 21554 399978
rect 21622 399922 21678 399978
rect 21250 382294 21306 382350
rect 21374 382294 21430 382350
rect 21498 382294 21554 382350
rect 21622 382294 21678 382350
rect 21250 382170 21306 382226
rect 21374 382170 21430 382226
rect 21498 382170 21554 382226
rect 21622 382170 21678 382226
rect 21250 382046 21306 382102
rect 21374 382046 21430 382102
rect 21498 382046 21554 382102
rect 21622 382046 21678 382102
rect 21250 381922 21306 381978
rect 21374 381922 21430 381978
rect 21498 381922 21554 381978
rect 21622 381922 21678 381978
rect 21250 364294 21306 364350
rect 21374 364294 21430 364350
rect 21498 364294 21554 364350
rect 21622 364294 21678 364350
rect 21250 364170 21306 364226
rect 21374 364170 21430 364226
rect 21498 364170 21554 364226
rect 21622 364170 21678 364226
rect 21250 364046 21306 364102
rect 21374 364046 21430 364102
rect 21498 364046 21554 364102
rect 21622 364046 21678 364102
rect 21250 363922 21306 363978
rect 21374 363922 21430 363978
rect 21498 363922 21554 363978
rect 21622 363922 21678 363978
rect 21250 346294 21306 346350
rect 21374 346294 21430 346350
rect 21498 346294 21554 346350
rect 21622 346294 21678 346350
rect 21250 346170 21306 346226
rect 21374 346170 21430 346226
rect 21498 346170 21554 346226
rect 21622 346170 21678 346226
rect 21250 346046 21306 346102
rect 21374 346046 21430 346102
rect 21498 346046 21554 346102
rect 21622 346046 21678 346102
rect 21250 345922 21306 345978
rect 21374 345922 21430 345978
rect 21498 345922 21554 345978
rect 21622 345922 21678 345978
rect 21250 328294 21306 328350
rect 21374 328294 21430 328350
rect 21498 328294 21554 328350
rect 21622 328294 21678 328350
rect 21250 328170 21306 328226
rect 21374 328170 21430 328226
rect 21498 328170 21554 328226
rect 21622 328170 21678 328226
rect 21250 328046 21306 328102
rect 21374 328046 21430 328102
rect 21498 328046 21554 328102
rect 21622 328046 21678 328102
rect 21250 327922 21306 327978
rect 21374 327922 21430 327978
rect 21498 327922 21554 327978
rect 21622 327922 21678 327978
rect 21250 310294 21306 310350
rect 21374 310294 21430 310350
rect 21498 310294 21554 310350
rect 21622 310294 21678 310350
rect 21250 310170 21306 310226
rect 21374 310170 21430 310226
rect 21498 310170 21554 310226
rect 21622 310170 21678 310226
rect 21250 310046 21306 310102
rect 21374 310046 21430 310102
rect 21498 310046 21554 310102
rect 21622 310046 21678 310102
rect 21250 309922 21306 309978
rect 21374 309922 21430 309978
rect 21498 309922 21554 309978
rect 21622 309922 21678 309978
rect 21250 292294 21306 292350
rect 21374 292294 21430 292350
rect 21498 292294 21554 292350
rect 21622 292294 21678 292350
rect 21250 292170 21306 292226
rect 21374 292170 21430 292226
rect 21498 292170 21554 292226
rect 21622 292170 21678 292226
rect 21250 292046 21306 292102
rect 21374 292046 21430 292102
rect 21498 292046 21554 292102
rect 21622 292046 21678 292102
rect 21250 291922 21306 291978
rect 21374 291922 21430 291978
rect 21498 291922 21554 291978
rect 21622 291922 21678 291978
rect 21250 274294 21306 274350
rect 21374 274294 21430 274350
rect 21498 274294 21554 274350
rect 21622 274294 21678 274350
rect 21250 274170 21306 274226
rect 21374 274170 21430 274226
rect 21498 274170 21554 274226
rect 21622 274170 21678 274226
rect 21250 274046 21306 274102
rect 21374 274046 21430 274102
rect 21498 274046 21554 274102
rect 21622 274046 21678 274102
rect 21250 273922 21306 273978
rect 21374 273922 21430 273978
rect 21498 273922 21554 273978
rect 21622 273922 21678 273978
rect 21250 256294 21306 256350
rect 21374 256294 21430 256350
rect 21498 256294 21554 256350
rect 21622 256294 21678 256350
rect 21250 256170 21306 256226
rect 21374 256170 21430 256226
rect 21498 256170 21554 256226
rect 21622 256170 21678 256226
rect 21250 256046 21306 256102
rect 21374 256046 21430 256102
rect 21498 256046 21554 256102
rect 21622 256046 21678 256102
rect 21250 255922 21306 255978
rect 21374 255922 21430 255978
rect 21498 255922 21554 255978
rect 21622 255922 21678 255978
rect 21250 238294 21306 238350
rect 21374 238294 21430 238350
rect 21498 238294 21554 238350
rect 21622 238294 21678 238350
rect 21250 238170 21306 238226
rect 21374 238170 21430 238226
rect 21498 238170 21554 238226
rect 21622 238170 21678 238226
rect 21250 238046 21306 238102
rect 21374 238046 21430 238102
rect 21498 238046 21554 238102
rect 21622 238046 21678 238102
rect 21250 237922 21306 237978
rect 21374 237922 21430 237978
rect 21498 237922 21554 237978
rect 21622 237922 21678 237978
rect 21250 220294 21306 220350
rect 21374 220294 21430 220350
rect 21498 220294 21554 220350
rect 21622 220294 21678 220350
rect 21250 220170 21306 220226
rect 21374 220170 21430 220226
rect 21498 220170 21554 220226
rect 21622 220170 21678 220226
rect 21250 220046 21306 220102
rect 21374 220046 21430 220102
rect 21498 220046 21554 220102
rect 21622 220046 21678 220102
rect 21250 219922 21306 219978
rect 21374 219922 21430 219978
rect 21498 219922 21554 219978
rect 21622 219922 21678 219978
rect 21250 202294 21306 202350
rect 21374 202294 21430 202350
rect 21498 202294 21554 202350
rect 21622 202294 21678 202350
rect 21250 202170 21306 202226
rect 21374 202170 21430 202226
rect 21498 202170 21554 202226
rect 21622 202170 21678 202226
rect 21250 202046 21306 202102
rect 21374 202046 21430 202102
rect 21498 202046 21554 202102
rect 21622 202046 21678 202102
rect 21250 201922 21306 201978
rect 21374 201922 21430 201978
rect 21498 201922 21554 201978
rect 21622 201922 21678 201978
rect 21250 184294 21306 184350
rect 21374 184294 21430 184350
rect 21498 184294 21554 184350
rect 21622 184294 21678 184350
rect 21250 184170 21306 184226
rect 21374 184170 21430 184226
rect 21498 184170 21554 184226
rect 21622 184170 21678 184226
rect 21250 184046 21306 184102
rect 21374 184046 21430 184102
rect 21498 184046 21554 184102
rect 21622 184046 21678 184102
rect 21250 183922 21306 183978
rect 21374 183922 21430 183978
rect 21498 183922 21554 183978
rect 21622 183922 21678 183978
rect 21250 166294 21306 166350
rect 21374 166294 21430 166350
rect 21498 166294 21554 166350
rect 21622 166294 21678 166350
rect 21250 166170 21306 166226
rect 21374 166170 21430 166226
rect 21498 166170 21554 166226
rect 21622 166170 21678 166226
rect 21250 166046 21306 166102
rect 21374 166046 21430 166102
rect 21498 166046 21554 166102
rect 21622 166046 21678 166102
rect 21250 165922 21306 165978
rect 21374 165922 21430 165978
rect 21498 165922 21554 165978
rect 21622 165922 21678 165978
rect 21250 148294 21306 148350
rect 21374 148294 21430 148350
rect 21498 148294 21554 148350
rect 21622 148294 21678 148350
rect 21250 148170 21306 148226
rect 21374 148170 21430 148226
rect 21498 148170 21554 148226
rect 21622 148170 21678 148226
rect 21250 148046 21306 148102
rect 21374 148046 21430 148102
rect 21498 148046 21554 148102
rect 21622 148046 21678 148102
rect 21250 147922 21306 147978
rect 21374 147922 21430 147978
rect 21498 147922 21554 147978
rect 21622 147922 21678 147978
rect 21250 130294 21306 130350
rect 21374 130294 21430 130350
rect 21498 130294 21554 130350
rect 21622 130294 21678 130350
rect 21250 130170 21306 130226
rect 21374 130170 21430 130226
rect 21498 130170 21554 130226
rect 21622 130170 21678 130226
rect 21250 130046 21306 130102
rect 21374 130046 21430 130102
rect 21498 130046 21554 130102
rect 21622 130046 21678 130102
rect 21250 129922 21306 129978
rect 21374 129922 21430 129978
rect 21498 129922 21554 129978
rect 21622 129922 21678 129978
rect 21250 112294 21306 112350
rect 21374 112294 21430 112350
rect 21498 112294 21554 112350
rect 21622 112294 21678 112350
rect 21250 112170 21306 112226
rect 21374 112170 21430 112226
rect 21498 112170 21554 112226
rect 21622 112170 21678 112226
rect 21250 112046 21306 112102
rect 21374 112046 21430 112102
rect 21498 112046 21554 112102
rect 21622 112046 21678 112102
rect 21250 111922 21306 111978
rect 21374 111922 21430 111978
rect 21498 111922 21554 111978
rect 21622 111922 21678 111978
rect 21250 94294 21306 94350
rect 21374 94294 21430 94350
rect 21498 94294 21554 94350
rect 21622 94294 21678 94350
rect 21250 94170 21306 94226
rect 21374 94170 21430 94226
rect 21498 94170 21554 94226
rect 21622 94170 21678 94226
rect 21250 94046 21306 94102
rect 21374 94046 21430 94102
rect 21498 94046 21554 94102
rect 21622 94046 21678 94102
rect 21250 93922 21306 93978
rect 21374 93922 21430 93978
rect 21498 93922 21554 93978
rect 21622 93922 21678 93978
rect 21250 76294 21306 76350
rect 21374 76294 21430 76350
rect 21498 76294 21554 76350
rect 21622 76294 21678 76350
rect 21250 76170 21306 76226
rect 21374 76170 21430 76226
rect 21498 76170 21554 76226
rect 21622 76170 21678 76226
rect 21250 76046 21306 76102
rect 21374 76046 21430 76102
rect 21498 76046 21554 76102
rect 21622 76046 21678 76102
rect 21250 75922 21306 75978
rect 21374 75922 21430 75978
rect 21498 75922 21554 75978
rect 21622 75922 21678 75978
rect 21250 58294 21306 58350
rect 21374 58294 21430 58350
rect 21498 58294 21554 58350
rect 21622 58294 21678 58350
rect 21250 58170 21306 58226
rect 21374 58170 21430 58226
rect 21498 58170 21554 58226
rect 21622 58170 21678 58226
rect 21250 58046 21306 58102
rect 21374 58046 21430 58102
rect 21498 58046 21554 58102
rect 21622 58046 21678 58102
rect 21250 57922 21306 57978
rect 21374 57922 21430 57978
rect 21498 57922 21554 57978
rect 21622 57922 21678 57978
rect 21250 40294 21306 40350
rect 21374 40294 21430 40350
rect 21498 40294 21554 40350
rect 21622 40294 21678 40350
rect 21250 40170 21306 40226
rect 21374 40170 21430 40226
rect 21498 40170 21554 40226
rect 21622 40170 21678 40226
rect 21250 40046 21306 40102
rect 21374 40046 21430 40102
rect 21498 40046 21554 40102
rect 21622 40046 21678 40102
rect 21250 39922 21306 39978
rect 21374 39922 21430 39978
rect 21498 39922 21554 39978
rect 21622 39922 21678 39978
rect 21250 22294 21306 22350
rect 21374 22294 21430 22350
rect 21498 22294 21554 22350
rect 21622 22294 21678 22350
rect 21250 22170 21306 22226
rect 21374 22170 21430 22226
rect 21498 22170 21554 22226
rect 21622 22170 21678 22226
rect 21250 22046 21306 22102
rect 21374 22046 21430 22102
rect 21498 22046 21554 22102
rect 21622 22046 21678 22102
rect 21250 21922 21306 21978
rect 21374 21922 21430 21978
rect 21498 21922 21554 21978
rect 21622 21922 21678 21978
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 24970 514294 25026 514350
rect 25094 514294 25150 514350
rect 25218 514294 25274 514350
rect 25342 514294 25398 514350
rect 24970 514170 25026 514226
rect 25094 514170 25150 514226
rect 25218 514170 25274 514226
rect 25342 514170 25398 514226
rect 24970 514046 25026 514102
rect 25094 514046 25150 514102
rect 25218 514046 25274 514102
rect 25342 514046 25398 514102
rect 24970 513922 25026 513978
rect 25094 513922 25150 513978
rect 25218 513922 25274 513978
rect 25342 513922 25398 513978
rect 24970 496294 25026 496350
rect 25094 496294 25150 496350
rect 25218 496294 25274 496350
rect 25342 496294 25398 496350
rect 24970 496170 25026 496226
rect 25094 496170 25150 496226
rect 25218 496170 25274 496226
rect 25342 496170 25398 496226
rect 24970 496046 25026 496102
rect 25094 496046 25150 496102
rect 25218 496046 25274 496102
rect 25342 496046 25398 496102
rect 24970 495922 25026 495978
rect 25094 495922 25150 495978
rect 25218 495922 25274 495978
rect 25342 495922 25398 495978
rect 24970 478294 25026 478350
rect 25094 478294 25150 478350
rect 25218 478294 25274 478350
rect 25342 478294 25398 478350
rect 24970 478170 25026 478226
rect 25094 478170 25150 478226
rect 25218 478170 25274 478226
rect 25342 478170 25398 478226
rect 24970 478046 25026 478102
rect 25094 478046 25150 478102
rect 25218 478046 25274 478102
rect 25342 478046 25398 478102
rect 24970 477922 25026 477978
rect 25094 477922 25150 477978
rect 25218 477922 25274 477978
rect 25342 477922 25398 477978
rect 24970 460294 25026 460350
rect 25094 460294 25150 460350
rect 25218 460294 25274 460350
rect 25342 460294 25398 460350
rect 24970 460170 25026 460226
rect 25094 460170 25150 460226
rect 25218 460170 25274 460226
rect 25342 460170 25398 460226
rect 24970 460046 25026 460102
rect 25094 460046 25150 460102
rect 25218 460046 25274 460102
rect 25342 460046 25398 460102
rect 24970 459922 25026 459978
rect 25094 459922 25150 459978
rect 25218 459922 25274 459978
rect 25342 459922 25398 459978
rect 24970 442294 25026 442350
rect 25094 442294 25150 442350
rect 25218 442294 25274 442350
rect 25342 442294 25398 442350
rect 24970 442170 25026 442226
rect 25094 442170 25150 442226
rect 25218 442170 25274 442226
rect 25342 442170 25398 442226
rect 24970 442046 25026 442102
rect 25094 442046 25150 442102
rect 25218 442046 25274 442102
rect 25342 442046 25398 442102
rect 24970 441922 25026 441978
rect 25094 441922 25150 441978
rect 25218 441922 25274 441978
rect 25342 441922 25398 441978
rect 24970 424294 25026 424350
rect 25094 424294 25150 424350
rect 25218 424294 25274 424350
rect 25342 424294 25398 424350
rect 24970 424170 25026 424226
rect 25094 424170 25150 424226
rect 25218 424170 25274 424226
rect 25342 424170 25398 424226
rect 24970 424046 25026 424102
rect 25094 424046 25150 424102
rect 25218 424046 25274 424102
rect 25342 424046 25398 424102
rect 24970 423922 25026 423978
rect 25094 423922 25150 423978
rect 25218 423922 25274 423978
rect 25342 423922 25398 423978
rect 24970 406294 25026 406350
rect 25094 406294 25150 406350
rect 25218 406294 25274 406350
rect 25342 406294 25398 406350
rect 24970 406170 25026 406226
rect 25094 406170 25150 406226
rect 25218 406170 25274 406226
rect 25342 406170 25398 406226
rect 24970 406046 25026 406102
rect 25094 406046 25150 406102
rect 25218 406046 25274 406102
rect 25342 406046 25398 406102
rect 24970 405922 25026 405978
rect 25094 405922 25150 405978
rect 25218 405922 25274 405978
rect 25342 405922 25398 405978
rect 24970 388294 25026 388350
rect 25094 388294 25150 388350
rect 25218 388294 25274 388350
rect 25342 388294 25398 388350
rect 24970 388170 25026 388226
rect 25094 388170 25150 388226
rect 25218 388170 25274 388226
rect 25342 388170 25398 388226
rect 24970 388046 25026 388102
rect 25094 388046 25150 388102
rect 25218 388046 25274 388102
rect 25342 388046 25398 388102
rect 24970 387922 25026 387978
rect 25094 387922 25150 387978
rect 25218 387922 25274 387978
rect 25342 387922 25398 387978
rect 24970 370294 25026 370350
rect 25094 370294 25150 370350
rect 25218 370294 25274 370350
rect 25342 370294 25398 370350
rect 24970 370170 25026 370226
rect 25094 370170 25150 370226
rect 25218 370170 25274 370226
rect 25342 370170 25398 370226
rect 24970 370046 25026 370102
rect 25094 370046 25150 370102
rect 25218 370046 25274 370102
rect 25342 370046 25398 370102
rect 24970 369922 25026 369978
rect 25094 369922 25150 369978
rect 25218 369922 25274 369978
rect 25342 369922 25398 369978
rect 24970 352294 25026 352350
rect 25094 352294 25150 352350
rect 25218 352294 25274 352350
rect 25342 352294 25398 352350
rect 24970 352170 25026 352226
rect 25094 352170 25150 352226
rect 25218 352170 25274 352226
rect 25342 352170 25398 352226
rect 24970 352046 25026 352102
rect 25094 352046 25150 352102
rect 25218 352046 25274 352102
rect 25342 352046 25398 352102
rect 24970 351922 25026 351978
rect 25094 351922 25150 351978
rect 25218 351922 25274 351978
rect 25342 351922 25398 351978
rect 24970 334294 25026 334350
rect 25094 334294 25150 334350
rect 25218 334294 25274 334350
rect 25342 334294 25398 334350
rect 24970 334170 25026 334226
rect 25094 334170 25150 334226
rect 25218 334170 25274 334226
rect 25342 334170 25398 334226
rect 24970 334046 25026 334102
rect 25094 334046 25150 334102
rect 25218 334046 25274 334102
rect 25342 334046 25398 334102
rect 24970 333922 25026 333978
rect 25094 333922 25150 333978
rect 25218 333922 25274 333978
rect 25342 333922 25398 333978
rect 24970 316294 25026 316350
rect 25094 316294 25150 316350
rect 25218 316294 25274 316350
rect 25342 316294 25398 316350
rect 24970 316170 25026 316226
rect 25094 316170 25150 316226
rect 25218 316170 25274 316226
rect 25342 316170 25398 316226
rect 24970 316046 25026 316102
rect 25094 316046 25150 316102
rect 25218 316046 25274 316102
rect 25342 316046 25398 316102
rect 24970 315922 25026 315978
rect 25094 315922 25150 315978
rect 25218 315922 25274 315978
rect 25342 315922 25398 315978
rect 24970 298294 25026 298350
rect 25094 298294 25150 298350
rect 25218 298294 25274 298350
rect 25342 298294 25398 298350
rect 24970 298170 25026 298226
rect 25094 298170 25150 298226
rect 25218 298170 25274 298226
rect 25342 298170 25398 298226
rect 24970 298046 25026 298102
rect 25094 298046 25150 298102
rect 25218 298046 25274 298102
rect 25342 298046 25398 298102
rect 24970 297922 25026 297978
rect 25094 297922 25150 297978
rect 25218 297922 25274 297978
rect 25342 297922 25398 297978
rect 24970 280294 25026 280350
rect 25094 280294 25150 280350
rect 25218 280294 25274 280350
rect 25342 280294 25398 280350
rect 24970 280170 25026 280226
rect 25094 280170 25150 280226
rect 25218 280170 25274 280226
rect 25342 280170 25398 280226
rect 24970 280046 25026 280102
rect 25094 280046 25150 280102
rect 25218 280046 25274 280102
rect 25342 280046 25398 280102
rect 24970 279922 25026 279978
rect 25094 279922 25150 279978
rect 25218 279922 25274 279978
rect 25342 279922 25398 279978
rect 24970 262294 25026 262350
rect 25094 262294 25150 262350
rect 25218 262294 25274 262350
rect 25342 262294 25398 262350
rect 24970 262170 25026 262226
rect 25094 262170 25150 262226
rect 25218 262170 25274 262226
rect 25342 262170 25398 262226
rect 24970 262046 25026 262102
rect 25094 262046 25150 262102
rect 25218 262046 25274 262102
rect 25342 262046 25398 262102
rect 24970 261922 25026 261978
rect 25094 261922 25150 261978
rect 25218 261922 25274 261978
rect 25342 261922 25398 261978
rect 24970 244294 25026 244350
rect 25094 244294 25150 244350
rect 25218 244294 25274 244350
rect 25342 244294 25398 244350
rect 24970 244170 25026 244226
rect 25094 244170 25150 244226
rect 25218 244170 25274 244226
rect 25342 244170 25398 244226
rect 24970 244046 25026 244102
rect 25094 244046 25150 244102
rect 25218 244046 25274 244102
rect 25342 244046 25398 244102
rect 24970 243922 25026 243978
rect 25094 243922 25150 243978
rect 25218 243922 25274 243978
rect 25342 243922 25398 243978
rect 24970 226294 25026 226350
rect 25094 226294 25150 226350
rect 25218 226294 25274 226350
rect 25342 226294 25398 226350
rect 24970 226170 25026 226226
rect 25094 226170 25150 226226
rect 25218 226170 25274 226226
rect 25342 226170 25398 226226
rect 24970 226046 25026 226102
rect 25094 226046 25150 226102
rect 25218 226046 25274 226102
rect 25342 226046 25398 226102
rect 24970 225922 25026 225978
rect 25094 225922 25150 225978
rect 25218 225922 25274 225978
rect 25342 225922 25398 225978
rect 24970 208294 25026 208350
rect 25094 208294 25150 208350
rect 25218 208294 25274 208350
rect 25342 208294 25398 208350
rect 24970 208170 25026 208226
rect 25094 208170 25150 208226
rect 25218 208170 25274 208226
rect 25342 208170 25398 208226
rect 24970 208046 25026 208102
rect 25094 208046 25150 208102
rect 25218 208046 25274 208102
rect 25342 208046 25398 208102
rect 24970 207922 25026 207978
rect 25094 207922 25150 207978
rect 25218 207922 25274 207978
rect 25342 207922 25398 207978
rect 24970 190294 25026 190350
rect 25094 190294 25150 190350
rect 25218 190294 25274 190350
rect 25342 190294 25398 190350
rect 24970 190170 25026 190226
rect 25094 190170 25150 190226
rect 25218 190170 25274 190226
rect 25342 190170 25398 190226
rect 24970 190046 25026 190102
rect 25094 190046 25150 190102
rect 25218 190046 25274 190102
rect 25342 190046 25398 190102
rect 24970 189922 25026 189978
rect 25094 189922 25150 189978
rect 25218 189922 25274 189978
rect 25342 189922 25398 189978
rect 24970 172294 25026 172350
rect 25094 172294 25150 172350
rect 25218 172294 25274 172350
rect 25342 172294 25398 172350
rect 24970 172170 25026 172226
rect 25094 172170 25150 172226
rect 25218 172170 25274 172226
rect 25342 172170 25398 172226
rect 24970 172046 25026 172102
rect 25094 172046 25150 172102
rect 25218 172046 25274 172102
rect 25342 172046 25398 172102
rect 24970 171922 25026 171978
rect 25094 171922 25150 171978
rect 25218 171922 25274 171978
rect 25342 171922 25398 171978
rect 24970 154294 25026 154350
rect 25094 154294 25150 154350
rect 25218 154294 25274 154350
rect 25342 154294 25398 154350
rect 24970 154170 25026 154226
rect 25094 154170 25150 154226
rect 25218 154170 25274 154226
rect 25342 154170 25398 154226
rect 24970 154046 25026 154102
rect 25094 154046 25150 154102
rect 25218 154046 25274 154102
rect 25342 154046 25398 154102
rect 24970 153922 25026 153978
rect 25094 153922 25150 153978
rect 25218 153922 25274 153978
rect 25342 153922 25398 153978
rect 24970 136294 25026 136350
rect 25094 136294 25150 136350
rect 25218 136294 25274 136350
rect 25342 136294 25398 136350
rect 24970 136170 25026 136226
rect 25094 136170 25150 136226
rect 25218 136170 25274 136226
rect 25342 136170 25398 136226
rect 24970 136046 25026 136102
rect 25094 136046 25150 136102
rect 25218 136046 25274 136102
rect 25342 136046 25398 136102
rect 24970 135922 25026 135978
rect 25094 135922 25150 135978
rect 25218 135922 25274 135978
rect 25342 135922 25398 135978
rect 24970 118294 25026 118350
rect 25094 118294 25150 118350
rect 25218 118294 25274 118350
rect 25342 118294 25398 118350
rect 24970 118170 25026 118226
rect 25094 118170 25150 118226
rect 25218 118170 25274 118226
rect 25342 118170 25398 118226
rect 24970 118046 25026 118102
rect 25094 118046 25150 118102
rect 25218 118046 25274 118102
rect 25342 118046 25398 118102
rect 24970 117922 25026 117978
rect 25094 117922 25150 117978
rect 25218 117922 25274 117978
rect 25342 117922 25398 117978
rect 24970 100294 25026 100350
rect 25094 100294 25150 100350
rect 25218 100294 25274 100350
rect 25342 100294 25398 100350
rect 24970 100170 25026 100226
rect 25094 100170 25150 100226
rect 25218 100170 25274 100226
rect 25342 100170 25398 100226
rect 24970 100046 25026 100102
rect 25094 100046 25150 100102
rect 25218 100046 25274 100102
rect 25342 100046 25398 100102
rect 24970 99922 25026 99978
rect 25094 99922 25150 99978
rect 25218 99922 25274 99978
rect 25342 99922 25398 99978
rect 24970 82294 25026 82350
rect 25094 82294 25150 82350
rect 25218 82294 25274 82350
rect 25342 82294 25398 82350
rect 24970 82170 25026 82226
rect 25094 82170 25150 82226
rect 25218 82170 25274 82226
rect 25342 82170 25398 82226
rect 24970 82046 25026 82102
rect 25094 82046 25150 82102
rect 25218 82046 25274 82102
rect 25342 82046 25398 82102
rect 24970 81922 25026 81978
rect 25094 81922 25150 81978
rect 25218 81922 25274 81978
rect 25342 81922 25398 81978
rect 24970 64294 25026 64350
rect 25094 64294 25150 64350
rect 25218 64294 25274 64350
rect 25342 64294 25398 64350
rect 24970 64170 25026 64226
rect 25094 64170 25150 64226
rect 25218 64170 25274 64226
rect 25342 64170 25398 64226
rect 24970 64046 25026 64102
rect 25094 64046 25150 64102
rect 25218 64046 25274 64102
rect 25342 64046 25398 64102
rect 24970 63922 25026 63978
rect 25094 63922 25150 63978
rect 25218 63922 25274 63978
rect 25342 63922 25398 63978
rect 24970 46294 25026 46350
rect 25094 46294 25150 46350
rect 25218 46294 25274 46350
rect 25342 46294 25398 46350
rect 24970 46170 25026 46226
rect 25094 46170 25150 46226
rect 25218 46170 25274 46226
rect 25342 46170 25398 46226
rect 24970 46046 25026 46102
rect 25094 46046 25150 46102
rect 25218 46046 25274 46102
rect 25342 46046 25398 46102
rect 24970 45922 25026 45978
rect 25094 45922 25150 45978
rect 25218 45922 25274 45978
rect 25342 45922 25398 45978
rect 24970 28294 25026 28350
rect 25094 28294 25150 28350
rect 25218 28294 25274 28350
rect 25342 28294 25398 28350
rect 24970 28170 25026 28226
rect 25094 28170 25150 28226
rect 25218 28170 25274 28226
rect 25342 28170 25398 28226
rect 24970 28046 25026 28102
rect 25094 28046 25150 28102
rect 25218 28046 25274 28102
rect 25342 28046 25398 28102
rect 24970 27922 25026 27978
rect 25094 27922 25150 27978
rect 25218 27922 25274 27978
rect 25342 27922 25398 27978
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 39250 508294 39306 508350
rect 39374 508294 39430 508350
rect 39498 508294 39554 508350
rect 39622 508294 39678 508350
rect 39250 508170 39306 508226
rect 39374 508170 39430 508226
rect 39498 508170 39554 508226
rect 39622 508170 39678 508226
rect 39250 508046 39306 508102
rect 39374 508046 39430 508102
rect 39498 508046 39554 508102
rect 39622 508046 39678 508102
rect 39250 507922 39306 507978
rect 39374 507922 39430 507978
rect 39498 507922 39554 507978
rect 39622 507922 39678 507978
rect 39250 490294 39306 490350
rect 39374 490294 39430 490350
rect 39498 490294 39554 490350
rect 39622 490294 39678 490350
rect 39250 490170 39306 490226
rect 39374 490170 39430 490226
rect 39498 490170 39554 490226
rect 39622 490170 39678 490226
rect 39250 490046 39306 490102
rect 39374 490046 39430 490102
rect 39498 490046 39554 490102
rect 39622 490046 39678 490102
rect 39250 489922 39306 489978
rect 39374 489922 39430 489978
rect 39498 489922 39554 489978
rect 39622 489922 39678 489978
rect 39250 472294 39306 472350
rect 39374 472294 39430 472350
rect 39498 472294 39554 472350
rect 39622 472294 39678 472350
rect 39250 472170 39306 472226
rect 39374 472170 39430 472226
rect 39498 472170 39554 472226
rect 39622 472170 39678 472226
rect 39250 472046 39306 472102
rect 39374 472046 39430 472102
rect 39498 472046 39554 472102
rect 39622 472046 39678 472102
rect 39250 471922 39306 471978
rect 39374 471922 39430 471978
rect 39498 471922 39554 471978
rect 39622 471922 39678 471978
rect 39250 454294 39306 454350
rect 39374 454294 39430 454350
rect 39498 454294 39554 454350
rect 39622 454294 39678 454350
rect 39250 454170 39306 454226
rect 39374 454170 39430 454226
rect 39498 454170 39554 454226
rect 39622 454170 39678 454226
rect 39250 454046 39306 454102
rect 39374 454046 39430 454102
rect 39498 454046 39554 454102
rect 39622 454046 39678 454102
rect 39250 453922 39306 453978
rect 39374 453922 39430 453978
rect 39498 453922 39554 453978
rect 39622 453922 39678 453978
rect 39250 436294 39306 436350
rect 39374 436294 39430 436350
rect 39498 436294 39554 436350
rect 39622 436294 39678 436350
rect 39250 436170 39306 436226
rect 39374 436170 39430 436226
rect 39498 436170 39554 436226
rect 39622 436170 39678 436226
rect 39250 436046 39306 436102
rect 39374 436046 39430 436102
rect 39498 436046 39554 436102
rect 39622 436046 39678 436102
rect 39250 435922 39306 435978
rect 39374 435922 39430 435978
rect 39498 435922 39554 435978
rect 39622 435922 39678 435978
rect 39250 418294 39306 418350
rect 39374 418294 39430 418350
rect 39498 418294 39554 418350
rect 39622 418294 39678 418350
rect 39250 418170 39306 418226
rect 39374 418170 39430 418226
rect 39498 418170 39554 418226
rect 39622 418170 39678 418226
rect 39250 418046 39306 418102
rect 39374 418046 39430 418102
rect 39498 418046 39554 418102
rect 39622 418046 39678 418102
rect 39250 417922 39306 417978
rect 39374 417922 39430 417978
rect 39498 417922 39554 417978
rect 39622 417922 39678 417978
rect 39250 400294 39306 400350
rect 39374 400294 39430 400350
rect 39498 400294 39554 400350
rect 39622 400294 39678 400350
rect 39250 400170 39306 400226
rect 39374 400170 39430 400226
rect 39498 400170 39554 400226
rect 39622 400170 39678 400226
rect 39250 400046 39306 400102
rect 39374 400046 39430 400102
rect 39498 400046 39554 400102
rect 39622 400046 39678 400102
rect 39250 399922 39306 399978
rect 39374 399922 39430 399978
rect 39498 399922 39554 399978
rect 39622 399922 39678 399978
rect 39250 382294 39306 382350
rect 39374 382294 39430 382350
rect 39498 382294 39554 382350
rect 39622 382294 39678 382350
rect 39250 382170 39306 382226
rect 39374 382170 39430 382226
rect 39498 382170 39554 382226
rect 39622 382170 39678 382226
rect 39250 382046 39306 382102
rect 39374 382046 39430 382102
rect 39498 382046 39554 382102
rect 39622 382046 39678 382102
rect 39250 381922 39306 381978
rect 39374 381922 39430 381978
rect 39498 381922 39554 381978
rect 39622 381922 39678 381978
rect 39250 364294 39306 364350
rect 39374 364294 39430 364350
rect 39498 364294 39554 364350
rect 39622 364294 39678 364350
rect 39250 364170 39306 364226
rect 39374 364170 39430 364226
rect 39498 364170 39554 364226
rect 39622 364170 39678 364226
rect 39250 364046 39306 364102
rect 39374 364046 39430 364102
rect 39498 364046 39554 364102
rect 39622 364046 39678 364102
rect 39250 363922 39306 363978
rect 39374 363922 39430 363978
rect 39498 363922 39554 363978
rect 39622 363922 39678 363978
rect 39250 346294 39306 346350
rect 39374 346294 39430 346350
rect 39498 346294 39554 346350
rect 39622 346294 39678 346350
rect 39250 346170 39306 346226
rect 39374 346170 39430 346226
rect 39498 346170 39554 346226
rect 39622 346170 39678 346226
rect 39250 346046 39306 346102
rect 39374 346046 39430 346102
rect 39498 346046 39554 346102
rect 39622 346046 39678 346102
rect 39250 345922 39306 345978
rect 39374 345922 39430 345978
rect 39498 345922 39554 345978
rect 39622 345922 39678 345978
rect 39250 328294 39306 328350
rect 39374 328294 39430 328350
rect 39498 328294 39554 328350
rect 39622 328294 39678 328350
rect 39250 328170 39306 328226
rect 39374 328170 39430 328226
rect 39498 328170 39554 328226
rect 39622 328170 39678 328226
rect 39250 328046 39306 328102
rect 39374 328046 39430 328102
rect 39498 328046 39554 328102
rect 39622 328046 39678 328102
rect 39250 327922 39306 327978
rect 39374 327922 39430 327978
rect 39498 327922 39554 327978
rect 39622 327922 39678 327978
rect 39250 310294 39306 310350
rect 39374 310294 39430 310350
rect 39498 310294 39554 310350
rect 39622 310294 39678 310350
rect 39250 310170 39306 310226
rect 39374 310170 39430 310226
rect 39498 310170 39554 310226
rect 39622 310170 39678 310226
rect 39250 310046 39306 310102
rect 39374 310046 39430 310102
rect 39498 310046 39554 310102
rect 39622 310046 39678 310102
rect 39250 309922 39306 309978
rect 39374 309922 39430 309978
rect 39498 309922 39554 309978
rect 39622 309922 39678 309978
rect 39250 292294 39306 292350
rect 39374 292294 39430 292350
rect 39498 292294 39554 292350
rect 39622 292294 39678 292350
rect 39250 292170 39306 292226
rect 39374 292170 39430 292226
rect 39498 292170 39554 292226
rect 39622 292170 39678 292226
rect 39250 292046 39306 292102
rect 39374 292046 39430 292102
rect 39498 292046 39554 292102
rect 39622 292046 39678 292102
rect 39250 291922 39306 291978
rect 39374 291922 39430 291978
rect 39498 291922 39554 291978
rect 39622 291922 39678 291978
rect 39250 274294 39306 274350
rect 39374 274294 39430 274350
rect 39498 274294 39554 274350
rect 39622 274294 39678 274350
rect 39250 274170 39306 274226
rect 39374 274170 39430 274226
rect 39498 274170 39554 274226
rect 39622 274170 39678 274226
rect 39250 274046 39306 274102
rect 39374 274046 39430 274102
rect 39498 274046 39554 274102
rect 39622 274046 39678 274102
rect 39250 273922 39306 273978
rect 39374 273922 39430 273978
rect 39498 273922 39554 273978
rect 39622 273922 39678 273978
rect 39250 256294 39306 256350
rect 39374 256294 39430 256350
rect 39498 256294 39554 256350
rect 39622 256294 39678 256350
rect 39250 256170 39306 256226
rect 39374 256170 39430 256226
rect 39498 256170 39554 256226
rect 39622 256170 39678 256226
rect 39250 256046 39306 256102
rect 39374 256046 39430 256102
rect 39498 256046 39554 256102
rect 39622 256046 39678 256102
rect 39250 255922 39306 255978
rect 39374 255922 39430 255978
rect 39498 255922 39554 255978
rect 39622 255922 39678 255978
rect 39250 238294 39306 238350
rect 39374 238294 39430 238350
rect 39498 238294 39554 238350
rect 39622 238294 39678 238350
rect 39250 238170 39306 238226
rect 39374 238170 39430 238226
rect 39498 238170 39554 238226
rect 39622 238170 39678 238226
rect 39250 238046 39306 238102
rect 39374 238046 39430 238102
rect 39498 238046 39554 238102
rect 39622 238046 39678 238102
rect 39250 237922 39306 237978
rect 39374 237922 39430 237978
rect 39498 237922 39554 237978
rect 39622 237922 39678 237978
rect 39250 220294 39306 220350
rect 39374 220294 39430 220350
rect 39498 220294 39554 220350
rect 39622 220294 39678 220350
rect 39250 220170 39306 220226
rect 39374 220170 39430 220226
rect 39498 220170 39554 220226
rect 39622 220170 39678 220226
rect 39250 220046 39306 220102
rect 39374 220046 39430 220102
rect 39498 220046 39554 220102
rect 39622 220046 39678 220102
rect 39250 219922 39306 219978
rect 39374 219922 39430 219978
rect 39498 219922 39554 219978
rect 39622 219922 39678 219978
rect 39250 202294 39306 202350
rect 39374 202294 39430 202350
rect 39498 202294 39554 202350
rect 39622 202294 39678 202350
rect 39250 202170 39306 202226
rect 39374 202170 39430 202226
rect 39498 202170 39554 202226
rect 39622 202170 39678 202226
rect 39250 202046 39306 202102
rect 39374 202046 39430 202102
rect 39498 202046 39554 202102
rect 39622 202046 39678 202102
rect 39250 201922 39306 201978
rect 39374 201922 39430 201978
rect 39498 201922 39554 201978
rect 39622 201922 39678 201978
rect 39250 184294 39306 184350
rect 39374 184294 39430 184350
rect 39498 184294 39554 184350
rect 39622 184294 39678 184350
rect 39250 184170 39306 184226
rect 39374 184170 39430 184226
rect 39498 184170 39554 184226
rect 39622 184170 39678 184226
rect 39250 184046 39306 184102
rect 39374 184046 39430 184102
rect 39498 184046 39554 184102
rect 39622 184046 39678 184102
rect 39250 183922 39306 183978
rect 39374 183922 39430 183978
rect 39498 183922 39554 183978
rect 39622 183922 39678 183978
rect 39250 166294 39306 166350
rect 39374 166294 39430 166350
rect 39498 166294 39554 166350
rect 39622 166294 39678 166350
rect 39250 166170 39306 166226
rect 39374 166170 39430 166226
rect 39498 166170 39554 166226
rect 39622 166170 39678 166226
rect 39250 166046 39306 166102
rect 39374 166046 39430 166102
rect 39498 166046 39554 166102
rect 39622 166046 39678 166102
rect 39250 165922 39306 165978
rect 39374 165922 39430 165978
rect 39498 165922 39554 165978
rect 39622 165922 39678 165978
rect 39250 148294 39306 148350
rect 39374 148294 39430 148350
rect 39498 148294 39554 148350
rect 39622 148294 39678 148350
rect 39250 148170 39306 148226
rect 39374 148170 39430 148226
rect 39498 148170 39554 148226
rect 39622 148170 39678 148226
rect 39250 148046 39306 148102
rect 39374 148046 39430 148102
rect 39498 148046 39554 148102
rect 39622 148046 39678 148102
rect 39250 147922 39306 147978
rect 39374 147922 39430 147978
rect 39498 147922 39554 147978
rect 39622 147922 39678 147978
rect 39250 130294 39306 130350
rect 39374 130294 39430 130350
rect 39498 130294 39554 130350
rect 39622 130294 39678 130350
rect 39250 130170 39306 130226
rect 39374 130170 39430 130226
rect 39498 130170 39554 130226
rect 39622 130170 39678 130226
rect 39250 130046 39306 130102
rect 39374 130046 39430 130102
rect 39498 130046 39554 130102
rect 39622 130046 39678 130102
rect 39250 129922 39306 129978
rect 39374 129922 39430 129978
rect 39498 129922 39554 129978
rect 39622 129922 39678 129978
rect 39250 112294 39306 112350
rect 39374 112294 39430 112350
rect 39498 112294 39554 112350
rect 39622 112294 39678 112350
rect 39250 112170 39306 112226
rect 39374 112170 39430 112226
rect 39498 112170 39554 112226
rect 39622 112170 39678 112226
rect 39250 112046 39306 112102
rect 39374 112046 39430 112102
rect 39498 112046 39554 112102
rect 39622 112046 39678 112102
rect 39250 111922 39306 111978
rect 39374 111922 39430 111978
rect 39498 111922 39554 111978
rect 39622 111922 39678 111978
rect 39250 94294 39306 94350
rect 39374 94294 39430 94350
rect 39498 94294 39554 94350
rect 39622 94294 39678 94350
rect 39250 94170 39306 94226
rect 39374 94170 39430 94226
rect 39498 94170 39554 94226
rect 39622 94170 39678 94226
rect 39250 94046 39306 94102
rect 39374 94046 39430 94102
rect 39498 94046 39554 94102
rect 39622 94046 39678 94102
rect 39250 93922 39306 93978
rect 39374 93922 39430 93978
rect 39498 93922 39554 93978
rect 39622 93922 39678 93978
rect 39250 76294 39306 76350
rect 39374 76294 39430 76350
rect 39498 76294 39554 76350
rect 39622 76294 39678 76350
rect 39250 76170 39306 76226
rect 39374 76170 39430 76226
rect 39498 76170 39554 76226
rect 39622 76170 39678 76226
rect 39250 76046 39306 76102
rect 39374 76046 39430 76102
rect 39498 76046 39554 76102
rect 39622 76046 39678 76102
rect 39250 75922 39306 75978
rect 39374 75922 39430 75978
rect 39498 75922 39554 75978
rect 39622 75922 39678 75978
rect 39250 58294 39306 58350
rect 39374 58294 39430 58350
rect 39498 58294 39554 58350
rect 39622 58294 39678 58350
rect 39250 58170 39306 58226
rect 39374 58170 39430 58226
rect 39498 58170 39554 58226
rect 39622 58170 39678 58226
rect 39250 58046 39306 58102
rect 39374 58046 39430 58102
rect 39498 58046 39554 58102
rect 39622 58046 39678 58102
rect 39250 57922 39306 57978
rect 39374 57922 39430 57978
rect 39498 57922 39554 57978
rect 39622 57922 39678 57978
rect 39250 40294 39306 40350
rect 39374 40294 39430 40350
rect 39498 40294 39554 40350
rect 39622 40294 39678 40350
rect 39250 40170 39306 40226
rect 39374 40170 39430 40226
rect 39498 40170 39554 40226
rect 39622 40170 39678 40226
rect 39250 40046 39306 40102
rect 39374 40046 39430 40102
rect 39498 40046 39554 40102
rect 39622 40046 39678 40102
rect 39250 39922 39306 39978
rect 39374 39922 39430 39978
rect 39498 39922 39554 39978
rect 39622 39922 39678 39978
rect 39250 22294 39306 22350
rect 39374 22294 39430 22350
rect 39498 22294 39554 22350
rect 39622 22294 39678 22350
rect 39250 22170 39306 22226
rect 39374 22170 39430 22226
rect 39498 22170 39554 22226
rect 39622 22170 39678 22226
rect 39250 22046 39306 22102
rect 39374 22046 39430 22102
rect 39498 22046 39554 22102
rect 39622 22046 39678 22102
rect 39250 21922 39306 21978
rect 39374 21922 39430 21978
rect 39498 21922 39554 21978
rect 39622 21922 39678 21978
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 42970 514294 43026 514350
rect 43094 514294 43150 514350
rect 43218 514294 43274 514350
rect 43342 514294 43398 514350
rect 42970 514170 43026 514226
rect 43094 514170 43150 514226
rect 43218 514170 43274 514226
rect 43342 514170 43398 514226
rect 42970 514046 43026 514102
rect 43094 514046 43150 514102
rect 43218 514046 43274 514102
rect 43342 514046 43398 514102
rect 42970 513922 43026 513978
rect 43094 513922 43150 513978
rect 43218 513922 43274 513978
rect 43342 513922 43398 513978
rect 42970 496294 43026 496350
rect 43094 496294 43150 496350
rect 43218 496294 43274 496350
rect 43342 496294 43398 496350
rect 42970 496170 43026 496226
rect 43094 496170 43150 496226
rect 43218 496170 43274 496226
rect 43342 496170 43398 496226
rect 42970 496046 43026 496102
rect 43094 496046 43150 496102
rect 43218 496046 43274 496102
rect 43342 496046 43398 496102
rect 42970 495922 43026 495978
rect 43094 495922 43150 495978
rect 43218 495922 43274 495978
rect 43342 495922 43398 495978
rect 42970 478294 43026 478350
rect 43094 478294 43150 478350
rect 43218 478294 43274 478350
rect 43342 478294 43398 478350
rect 42970 478170 43026 478226
rect 43094 478170 43150 478226
rect 43218 478170 43274 478226
rect 43342 478170 43398 478226
rect 42970 478046 43026 478102
rect 43094 478046 43150 478102
rect 43218 478046 43274 478102
rect 43342 478046 43398 478102
rect 42970 477922 43026 477978
rect 43094 477922 43150 477978
rect 43218 477922 43274 477978
rect 43342 477922 43398 477978
rect 42970 460294 43026 460350
rect 43094 460294 43150 460350
rect 43218 460294 43274 460350
rect 43342 460294 43398 460350
rect 42970 460170 43026 460226
rect 43094 460170 43150 460226
rect 43218 460170 43274 460226
rect 43342 460170 43398 460226
rect 42970 460046 43026 460102
rect 43094 460046 43150 460102
rect 43218 460046 43274 460102
rect 43342 460046 43398 460102
rect 42970 459922 43026 459978
rect 43094 459922 43150 459978
rect 43218 459922 43274 459978
rect 43342 459922 43398 459978
rect 42970 442294 43026 442350
rect 43094 442294 43150 442350
rect 43218 442294 43274 442350
rect 43342 442294 43398 442350
rect 42970 442170 43026 442226
rect 43094 442170 43150 442226
rect 43218 442170 43274 442226
rect 43342 442170 43398 442226
rect 42970 442046 43026 442102
rect 43094 442046 43150 442102
rect 43218 442046 43274 442102
rect 43342 442046 43398 442102
rect 42970 441922 43026 441978
rect 43094 441922 43150 441978
rect 43218 441922 43274 441978
rect 43342 441922 43398 441978
rect 42970 424294 43026 424350
rect 43094 424294 43150 424350
rect 43218 424294 43274 424350
rect 43342 424294 43398 424350
rect 42970 424170 43026 424226
rect 43094 424170 43150 424226
rect 43218 424170 43274 424226
rect 43342 424170 43398 424226
rect 42970 424046 43026 424102
rect 43094 424046 43150 424102
rect 43218 424046 43274 424102
rect 43342 424046 43398 424102
rect 42970 423922 43026 423978
rect 43094 423922 43150 423978
rect 43218 423922 43274 423978
rect 43342 423922 43398 423978
rect 42970 406294 43026 406350
rect 43094 406294 43150 406350
rect 43218 406294 43274 406350
rect 43342 406294 43398 406350
rect 42970 406170 43026 406226
rect 43094 406170 43150 406226
rect 43218 406170 43274 406226
rect 43342 406170 43398 406226
rect 42970 406046 43026 406102
rect 43094 406046 43150 406102
rect 43218 406046 43274 406102
rect 43342 406046 43398 406102
rect 42970 405922 43026 405978
rect 43094 405922 43150 405978
rect 43218 405922 43274 405978
rect 43342 405922 43398 405978
rect 42970 388294 43026 388350
rect 43094 388294 43150 388350
rect 43218 388294 43274 388350
rect 43342 388294 43398 388350
rect 42970 388170 43026 388226
rect 43094 388170 43150 388226
rect 43218 388170 43274 388226
rect 43342 388170 43398 388226
rect 42970 388046 43026 388102
rect 43094 388046 43150 388102
rect 43218 388046 43274 388102
rect 43342 388046 43398 388102
rect 42970 387922 43026 387978
rect 43094 387922 43150 387978
rect 43218 387922 43274 387978
rect 43342 387922 43398 387978
rect 42970 370294 43026 370350
rect 43094 370294 43150 370350
rect 43218 370294 43274 370350
rect 43342 370294 43398 370350
rect 42970 370170 43026 370226
rect 43094 370170 43150 370226
rect 43218 370170 43274 370226
rect 43342 370170 43398 370226
rect 42970 370046 43026 370102
rect 43094 370046 43150 370102
rect 43218 370046 43274 370102
rect 43342 370046 43398 370102
rect 42970 369922 43026 369978
rect 43094 369922 43150 369978
rect 43218 369922 43274 369978
rect 43342 369922 43398 369978
rect 42970 352294 43026 352350
rect 43094 352294 43150 352350
rect 43218 352294 43274 352350
rect 43342 352294 43398 352350
rect 42970 352170 43026 352226
rect 43094 352170 43150 352226
rect 43218 352170 43274 352226
rect 43342 352170 43398 352226
rect 42970 352046 43026 352102
rect 43094 352046 43150 352102
rect 43218 352046 43274 352102
rect 43342 352046 43398 352102
rect 42970 351922 43026 351978
rect 43094 351922 43150 351978
rect 43218 351922 43274 351978
rect 43342 351922 43398 351978
rect 42970 334294 43026 334350
rect 43094 334294 43150 334350
rect 43218 334294 43274 334350
rect 43342 334294 43398 334350
rect 42970 334170 43026 334226
rect 43094 334170 43150 334226
rect 43218 334170 43274 334226
rect 43342 334170 43398 334226
rect 42970 334046 43026 334102
rect 43094 334046 43150 334102
rect 43218 334046 43274 334102
rect 43342 334046 43398 334102
rect 42970 333922 43026 333978
rect 43094 333922 43150 333978
rect 43218 333922 43274 333978
rect 43342 333922 43398 333978
rect 42970 316294 43026 316350
rect 43094 316294 43150 316350
rect 43218 316294 43274 316350
rect 43342 316294 43398 316350
rect 42970 316170 43026 316226
rect 43094 316170 43150 316226
rect 43218 316170 43274 316226
rect 43342 316170 43398 316226
rect 42970 316046 43026 316102
rect 43094 316046 43150 316102
rect 43218 316046 43274 316102
rect 43342 316046 43398 316102
rect 42970 315922 43026 315978
rect 43094 315922 43150 315978
rect 43218 315922 43274 315978
rect 43342 315922 43398 315978
rect 42970 298294 43026 298350
rect 43094 298294 43150 298350
rect 43218 298294 43274 298350
rect 43342 298294 43398 298350
rect 42970 298170 43026 298226
rect 43094 298170 43150 298226
rect 43218 298170 43274 298226
rect 43342 298170 43398 298226
rect 42970 298046 43026 298102
rect 43094 298046 43150 298102
rect 43218 298046 43274 298102
rect 43342 298046 43398 298102
rect 42970 297922 43026 297978
rect 43094 297922 43150 297978
rect 43218 297922 43274 297978
rect 43342 297922 43398 297978
rect 42970 280294 43026 280350
rect 43094 280294 43150 280350
rect 43218 280294 43274 280350
rect 43342 280294 43398 280350
rect 42970 280170 43026 280226
rect 43094 280170 43150 280226
rect 43218 280170 43274 280226
rect 43342 280170 43398 280226
rect 42970 280046 43026 280102
rect 43094 280046 43150 280102
rect 43218 280046 43274 280102
rect 43342 280046 43398 280102
rect 42970 279922 43026 279978
rect 43094 279922 43150 279978
rect 43218 279922 43274 279978
rect 43342 279922 43398 279978
rect 42970 262294 43026 262350
rect 43094 262294 43150 262350
rect 43218 262294 43274 262350
rect 43342 262294 43398 262350
rect 42970 262170 43026 262226
rect 43094 262170 43150 262226
rect 43218 262170 43274 262226
rect 43342 262170 43398 262226
rect 42970 262046 43026 262102
rect 43094 262046 43150 262102
rect 43218 262046 43274 262102
rect 43342 262046 43398 262102
rect 42970 261922 43026 261978
rect 43094 261922 43150 261978
rect 43218 261922 43274 261978
rect 43342 261922 43398 261978
rect 42970 244294 43026 244350
rect 43094 244294 43150 244350
rect 43218 244294 43274 244350
rect 43342 244294 43398 244350
rect 42970 244170 43026 244226
rect 43094 244170 43150 244226
rect 43218 244170 43274 244226
rect 43342 244170 43398 244226
rect 42970 244046 43026 244102
rect 43094 244046 43150 244102
rect 43218 244046 43274 244102
rect 43342 244046 43398 244102
rect 42970 243922 43026 243978
rect 43094 243922 43150 243978
rect 43218 243922 43274 243978
rect 43342 243922 43398 243978
rect 42970 226294 43026 226350
rect 43094 226294 43150 226350
rect 43218 226294 43274 226350
rect 43342 226294 43398 226350
rect 42970 226170 43026 226226
rect 43094 226170 43150 226226
rect 43218 226170 43274 226226
rect 43342 226170 43398 226226
rect 42970 226046 43026 226102
rect 43094 226046 43150 226102
rect 43218 226046 43274 226102
rect 43342 226046 43398 226102
rect 42970 225922 43026 225978
rect 43094 225922 43150 225978
rect 43218 225922 43274 225978
rect 43342 225922 43398 225978
rect 42970 208294 43026 208350
rect 43094 208294 43150 208350
rect 43218 208294 43274 208350
rect 43342 208294 43398 208350
rect 42970 208170 43026 208226
rect 43094 208170 43150 208226
rect 43218 208170 43274 208226
rect 43342 208170 43398 208226
rect 42970 208046 43026 208102
rect 43094 208046 43150 208102
rect 43218 208046 43274 208102
rect 43342 208046 43398 208102
rect 42970 207922 43026 207978
rect 43094 207922 43150 207978
rect 43218 207922 43274 207978
rect 43342 207922 43398 207978
rect 42970 190294 43026 190350
rect 43094 190294 43150 190350
rect 43218 190294 43274 190350
rect 43342 190294 43398 190350
rect 42970 190170 43026 190226
rect 43094 190170 43150 190226
rect 43218 190170 43274 190226
rect 43342 190170 43398 190226
rect 42970 190046 43026 190102
rect 43094 190046 43150 190102
rect 43218 190046 43274 190102
rect 43342 190046 43398 190102
rect 42970 189922 43026 189978
rect 43094 189922 43150 189978
rect 43218 189922 43274 189978
rect 43342 189922 43398 189978
rect 42970 172294 43026 172350
rect 43094 172294 43150 172350
rect 43218 172294 43274 172350
rect 43342 172294 43398 172350
rect 42970 172170 43026 172226
rect 43094 172170 43150 172226
rect 43218 172170 43274 172226
rect 43342 172170 43398 172226
rect 42970 172046 43026 172102
rect 43094 172046 43150 172102
rect 43218 172046 43274 172102
rect 43342 172046 43398 172102
rect 42970 171922 43026 171978
rect 43094 171922 43150 171978
rect 43218 171922 43274 171978
rect 43342 171922 43398 171978
rect 42970 154294 43026 154350
rect 43094 154294 43150 154350
rect 43218 154294 43274 154350
rect 43342 154294 43398 154350
rect 42970 154170 43026 154226
rect 43094 154170 43150 154226
rect 43218 154170 43274 154226
rect 43342 154170 43398 154226
rect 42970 154046 43026 154102
rect 43094 154046 43150 154102
rect 43218 154046 43274 154102
rect 43342 154046 43398 154102
rect 42970 153922 43026 153978
rect 43094 153922 43150 153978
rect 43218 153922 43274 153978
rect 43342 153922 43398 153978
rect 42970 136294 43026 136350
rect 43094 136294 43150 136350
rect 43218 136294 43274 136350
rect 43342 136294 43398 136350
rect 42970 136170 43026 136226
rect 43094 136170 43150 136226
rect 43218 136170 43274 136226
rect 43342 136170 43398 136226
rect 42970 136046 43026 136102
rect 43094 136046 43150 136102
rect 43218 136046 43274 136102
rect 43342 136046 43398 136102
rect 42970 135922 43026 135978
rect 43094 135922 43150 135978
rect 43218 135922 43274 135978
rect 43342 135922 43398 135978
rect 42970 118294 43026 118350
rect 43094 118294 43150 118350
rect 43218 118294 43274 118350
rect 43342 118294 43398 118350
rect 42970 118170 43026 118226
rect 43094 118170 43150 118226
rect 43218 118170 43274 118226
rect 43342 118170 43398 118226
rect 42970 118046 43026 118102
rect 43094 118046 43150 118102
rect 43218 118046 43274 118102
rect 43342 118046 43398 118102
rect 42970 117922 43026 117978
rect 43094 117922 43150 117978
rect 43218 117922 43274 117978
rect 43342 117922 43398 117978
rect 42970 100294 43026 100350
rect 43094 100294 43150 100350
rect 43218 100294 43274 100350
rect 43342 100294 43398 100350
rect 42970 100170 43026 100226
rect 43094 100170 43150 100226
rect 43218 100170 43274 100226
rect 43342 100170 43398 100226
rect 42970 100046 43026 100102
rect 43094 100046 43150 100102
rect 43218 100046 43274 100102
rect 43342 100046 43398 100102
rect 42970 99922 43026 99978
rect 43094 99922 43150 99978
rect 43218 99922 43274 99978
rect 43342 99922 43398 99978
rect 42970 82294 43026 82350
rect 43094 82294 43150 82350
rect 43218 82294 43274 82350
rect 43342 82294 43398 82350
rect 42970 82170 43026 82226
rect 43094 82170 43150 82226
rect 43218 82170 43274 82226
rect 43342 82170 43398 82226
rect 42970 82046 43026 82102
rect 43094 82046 43150 82102
rect 43218 82046 43274 82102
rect 43342 82046 43398 82102
rect 42970 81922 43026 81978
rect 43094 81922 43150 81978
rect 43218 81922 43274 81978
rect 43342 81922 43398 81978
rect 42970 64294 43026 64350
rect 43094 64294 43150 64350
rect 43218 64294 43274 64350
rect 43342 64294 43398 64350
rect 42970 64170 43026 64226
rect 43094 64170 43150 64226
rect 43218 64170 43274 64226
rect 43342 64170 43398 64226
rect 42970 64046 43026 64102
rect 43094 64046 43150 64102
rect 43218 64046 43274 64102
rect 43342 64046 43398 64102
rect 42970 63922 43026 63978
rect 43094 63922 43150 63978
rect 43218 63922 43274 63978
rect 43342 63922 43398 63978
rect 42970 46294 43026 46350
rect 43094 46294 43150 46350
rect 43218 46294 43274 46350
rect 43342 46294 43398 46350
rect 42970 46170 43026 46226
rect 43094 46170 43150 46226
rect 43218 46170 43274 46226
rect 43342 46170 43398 46226
rect 42970 46046 43026 46102
rect 43094 46046 43150 46102
rect 43218 46046 43274 46102
rect 43342 46046 43398 46102
rect 42970 45922 43026 45978
rect 43094 45922 43150 45978
rect 43218 45922 43274 45978
rect 43342 45922 43398 45978
rect 42970 28294 43026 28350
rect 43094 28294 43150 28350
rect 43218 28294 43274 28350
rect 43342 28294 43398 28350
rect 42970 28170 43026 28226
rect 43094 28170 43150 28226
rect 43218 28170 43274 28226
rect 43342 28170 43398 28226
rect 42970 28046 43026 28102
rect 43094 28046 43150 28102
rect 43218 28046 43274 28102
rect 43342 28046 43398 28102
rect 42970 27922 43026 27978
rect 43094 27922 43150 27978
rect 43218 27922 43274 27978
rect 43342 27922 43398 27978
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 57250 508294 57306 508350
rect 57374 508294 57430 508350
rect 57498 508294 57554 508350
rect 57622 508294 57678 508350
rect 57250 508170 57306 508226
rect 57374 508170 57430 508226
rect 57498 508170 57554 508226
rect 57622 508170 57678 508226
rect 57250 508046 57306 508102
rect 57374 508046 57430 508102
rect 57498 508046 57554 508102
rect 57622 508046 57678 508102
rect 57250 507922 57306 507978
rect 57374 507922 57430 507978
rect 57498 507922 57554 507978
rect 57622 507922 57678 507978
rect 57250 490294 57306 490350
rect 57374 490294 57430 490350
rect 57498 490294 57554 490350
rect 57622 490294 57678 490350
rect 57250 490170 57306 490226
rect 57374 490170 57430 490226
rect 57498 490170 57554 490226
rect 57622 490170 57678 490226
rect 57250 490046 57306 490102
rect 57374 490046 57430 490102
rect 57498 490046 57554 490102
rect 57622 490046 57678 490102
rect 57250 489922 57306 489978
rect 57374 489922 57430 489978
rect 57498 489922 57554 489978
rect 57622 489922 57678 489978
rect 57250 472294 57306 472350
rect 57374 472294 57430 472350
rect 57498 472294 57554 472350
rect 57622 472294 57678 472350
rect 57250 472170 57306 472226
rect 57374 472170 57430 472226
rect 57498 472170 57554 472226
rect 57622 472170 57678 472226
rect 57250 472046 57306 472102
rect 57374 472046 57430 472102
rect 57498 472046 57554 472102
rect 57622 472046 57678 472102
rect 57250 471922 57306 471978
rect 57374 471922 57430 471978
rect 57498 471922 57554 471978
rect 57622 471922 57678 471978
rect 57250 454294 57306 454350
rect 57374 454294 57430 454350
rect 57498 454294 57554 454350
rect 57622 454294 57678 454350
rect 57250 454170 57306 454226
rect 57374 454170 57430 454226
rect 57498 454170 57554 454226
rect 57622 454170 57678 454226
rect 57250 454046 57306 454102
rect 57374 454046 57430 454102
rect 57498 454046 57554 454102
rect 57622 454046 57678 454102
rect 57250 453922 57306 453978
rect 57374 453922 57430 453978
rect 57498 453922 57554 453978
rect 57622 453922 57678 453978
rect 57250 436294 57306 436350
rect 57374 436294 57430 436350
rect 57498 436294 57554 436350
rect 57622 436294 57678 436350
rect 57250 436170 57306 436226
rect 57374 436170 57430 436226
rect 57498 436170 57554 436226
rect 57622 436170 57678 436226
rect 57250 436046 57306 436102
rect 57374 436046 57430 436102
rect 57498 436046 57554 436102
rect 57622 436046 57678 436102
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 60970 514294 61026 514350
rect 61094 514294 61150 514350
rect 61218 514294 61274 514350
rect 61342 514294 61398 514350
rect 60970 514170 61026 514226
rect 61094 514170 61150 514226
rect 61218 514170 61274 514226
rect 61342 514170 61398 514226
rect 60970 514046 61026 514102
rect 61094 514046 61150 514102
rect 61218 514046 61274 514102
rect 61342 514046 61398 514102
rect 60970 513922 61026 513978
rect 61094 513922 61150 513978
rect 61218 513922 61274 513978
rect 61342 513922 61398 513978
rect 60970 496294 61026 496350
rect 61094 496294 61150 496350
rect 61218 496294 61274 496350
rect 61342 496294 61398 496350
rect 60970 496170 61026 496226
rect 61094 496170 61150 496226
rect 61218 496170 61274 496226
rect 61342 496170 61398 496226
rect 60970 496046 61026 496102
rect 61094 496046 61150 496102
rect 61218 496046 61274 496102
rect 61342 496046 61398 496102
rect 60970 495922 61026 495978
rect 61094 495922 61150 495978
rect 61218 495922 61274 495978
rect 61342 495922 61398 495978
rect 60970 478294 61026 478350
rect 61094 478294 61150 478350
rect 61218 478294 61274 478350
rect 61342 478294 61398 478350
rect 60970 478170 61026 478226
rect 61094 478170 61150 478226
rect 61218 478170 61274 478226
rect 61342 478170 61398 478226
rect 60970 478046 61026 478102
rect 61094 478046 61150 478102
rect 61218 478046 61274 478102
rect 61342 478046 61398 478102
rect 60970 477922 61026 477978
rect 61094 477922 61150 477978
rect 61218 477922 61274 477978
rect 61342 477922 61398 477978
rect 60970 460294 61026 460350
rect 61094 460294 61150 460350
rect 61218 460294 61274 460350
rect 61342 460294 61398 460350
rect 60970 460170 61026 460226
rect 61094 460170 61150 460226
rect 61218 460170 61274 460226
rect 61342 460170 61398 460226
rect 60970 460046 61026 460102
rect 61094 460046 61150 460102
rect 61218 460046 61274 460102
rect 61342 460046 61398 460102
rect 60970 459922 61026 459978
rect 61094 459922 61150 459978
rect 61218 459922 61274 459978
rect 61342 459922 61398 459978
rect 60970 442294 61026 442350
rect 61094 442294 61150 442350
rect 61218 442294 61274 442350
rect 61342 442294 61398 442350
rect 60970 442170 61026 442226
rect 61094 442170 61150 442226
rect 61218 442170 61274 442226
rect 61342 442170 61398 442226
rect 60970 442046 61026 442102
rect 61094 442046 61150 442102
rect 61218 442046 61274 442102
rect 61342 442046 61398 442102
rect 60970 441922 61026 441978
rect 61094 441922 61150 441978
rect 61218 441922 61274 441978
rect 61342 441922 61398 441978
rect 75250 597156 75306 597212
rect 75374 597156 75430 597212
rect 75498 597156 75554 597212
rect 75622 597156 75678 597212
rect 75250 597032 75306 597088
rect 75374 597032 75430 597088
rect 75498 597032 75554 597088
rect 75622 597032 75678 597088
rect 75250 596908 75306 596964
rect 75374 596908 75430 596964
rect 75498 596908 75554 596964
rect 75622 596908 75678 596964
rect 75250 596784 75306 596840
rect 75374 596784 75430 596840
rect 75498 596784 75554 596840
rect 75622 596784 75678 596840
rect 75250 580294 75306 580350
rect 75374 580294 75430 580350
rect 75498 580294 75554 580350
rect 75622 580294 75678 580350
rect 75250 580170 75306 580226
rect 75374 580170 75430 580226
rect 75498 580170 75554 580226
rect 75622 580170 75678 580226
rect 75250 580046 75306 580102
rect 75374 580046 75430 580102
rect 75498 580046 75554 580102
rect 75622 580046 75678 580102
rect 75250 579922 75306 579978
rect 75374 579922 75430 579978
rect 75498 579922 75554 579978
rect 75622 579922 75678 579978
rect 75250 562294 75306 562350
rect 75374 562294 75430 562350
rect 75498 562294 75554 562350
rect 75622 562294 75678 562350
rect 75250 562170 75306 562226
rect 75374 562170 75430 562226
rect 75498 562170 75554 562226
rect 75622 562170 75678 562226
rect 75250 562046 75306 562102
rect 75374 562046 75430 562102
rect 75498 562046 75554 562102
rect 75622 562046 75678 562102
rect 75250 561922 75306 561978
rect 75374 561922 75430 561978
rect 75498 561922 75554 561978
rect 75622 561922 75678 561978
rect 75250 544294 75306 544350
rect 75374 544294 75430 544350
rect 75498 544294 75554 544350
rect 75622 544294 75678 544350
rect 75250 544170 75306 544226
rect 75374 544170 75430 544226
rect 75498 544170 75554 544226
rect 75622 544170 75678 544226
rect 75250 544046 75306 544102
rect 75374 544046 75430 544102
rect 75498 544046 75554 544102
rect 75622 544046 75678 544102
rect 75250 543922 75306 543978
rect 75374 543922 75430 543978
rect 75498 543922 75554 543978
rect 75622 543922 75678 543978
rect 75250 526294 75306 526350
rect 75374 526294 75430 526350
rect 75498 526294 75554 526350
rect 75622 526294 75678 526350
rect 75250 526170 75306 526226
rect 75374 526170 75430 526226
rect 75498 526170 75554 526226
rect 75622 526170 75678 526226
rect 75250 526046 75306 526102
rect 75374 526046 75430 526102
rect 75498 526046 75554 526102
rect 75622 526046 75678 526102
rect 75250 525922 75306 525978
rect 75374 525922 75430 525978
rect 75498 525922 75554 525978
rect 75622 525922 75678 525978
rect 75250 508294 75306 508350
rect 75374 508294 75430 508350
rect 75498 508294 75554 508350
rect 75622 508294 75678 508350
rect 75250 508170 75306 508226
rect 75374 508170 75430 508226
rect 75498 508170 75554 508226
rect 75622 508170 75678 508226
rect 75250 508046 75306 508102
rect 75374 508046 75430 508102
rect 75498 508046 75554 508102
rect 75622 508046 75678 508102
rect 75250 507922 75306 507978
rect 75374 507922 75430 507978
rect 75498 507922 75554 507978
rect 75622 507922 75678 507978
rect 75250 490294 75306 490350
rect 75374 490294 75430 490350
rect 75498 490294 75554 490350
rect 75622 490294 75678 490350
rect 75250 490170 75306 490226
rect 75374 490170 75430 490226
rect 75498 490170 75554 490226
rect 75622 490170 75678 490226
rect 75250 490046 75306 490102
rect 75374 490046 75430 490102
rect 75498 490046 75554 490102
rect 75622 490046 75678 490102
rect 75250 489922 75306 489978
rect 75374 489922 75430 489978
rect 75498 489922 75554 489978
rect 75622 489922 75678 489978
rect 75250 472294 75306 472350
rect 75374 472294 75430 472350
rect 75498 472294 75554 472350
rect 75622 472294 75678 472350
rect 75250 472170 75306 472226
rect 75374 472170 75430 472226
rect 75498 472170 75554 472226
rect 75622 472170 75678 472226
rect 75250 472046 75306 472102
rect 75374 472046 75430 472102
rect 75498 472046 75554 472102
rect 75622 472046 75678 472102
rect 75250 471922 75306 471978
rect 75374 471922 75430 471978
rect 75498 471922 75554 471978
rect 75622 471922 75678 471978
rect 75250 454294 75306 454350
rect 75374 454294 75430 454350
rect 75498 454294 75554 454350
rect 75622 454294 75678 454350
rect 75250 454170 75306 454226
rect 75374 454170 75430 454226
rect 75498 454170 75554 454226
rect 75622 454170 75678 454226
rect 75250 454046 75306 454102
rect 75374 454046 75430 454102
rect 75498 454046 75554 454102
rect 75622 454046 75678 454102
rect 75250 453922 75306 453978
rect 75374 453922 75430 453978
rect 75498 453922 75554 453978
rect 75622 453922 75678 453978
rect 64518 436261 64574 436317
rect 64642 436261 64698 436317
rect 64518 436137 64574 436193
rect 64642 436137 64698 436193
rect 64518 436013 64574 436069
rect 64642 436013 64698 436069
rect 57250 435922 57306 435978
rect 57374 435922 57430 435978
rect 57498 435922 57554 435978
rect 57622 435922 57678 435978
rect 75250 436322 75306 436378
rect 75374 436322 75430 436378
rect 75498 436322 75554 436378
rect 75622 436322 75678 436378
rect 75250 436198 75306 436254
rect 75374 436198 75430 436254
rect 75498 436198 75554 436254
rect 75622 436198 75678 436254
rect 75250 436074 75306 436130
rect 75374 436074 75430 436130
rect 75498 436074 75554 436130
rect 75622 436074 75678 436130
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 78970 514294 79026 514350
rect 79094 514294 79150 514350
rect 79218 514294 79274 514350
rect 79342 514294 79398 514350
rect 78970 514170 79026 514226
rect 79094 514170 79150 514226
rect 79218 514170 79274 514226
rect 79342 514170 79398 514226
rect 78970 514046 79026 514102
rect 79094 514046 79150 514102
rect 79218 514046 79274 514102
rect 79342 514046 79398 514102
rect 78970 513922 79026 513978
rect 79094 513922 79150 513978
rect 79218 513922 79274 513978
rect 79342 513922 79398 513978
rect 78970 496294 79026 496350
rect 79094 496294 79150 496350
rect 79218 496294 79274 496350
rect 79342 496294 79398 496350
rect 78970 496170 79026 496226
rect 79094 496170 79150 496226
rect 79218 496170 79274 496226
rect 79342 496170 79398 496226
rect 78970 496046 79026 496102
rect 79094 496046 79150 496102
rect 79218 496046 79274 496102
rect 79342 496046 79398 496102
rect 78970 495922 79026 495978
rect 79094 495922 79150 495978
rect 79218 495922 79274 495978
rect 79342 495922 79398 495978
rect 78970 478294 79026 478350
rect 79094 478294 79150 478350
rect 79218 478294 79274 478350
rect 79342 478294 79398 478350
rect 78970 478170 79026 478226
rect 79094 478170 79150 478226
rect 79218 478170 79274 478226
rect 79342 478170 79398 478226
rect 78970 478046 79026 478102
rect 79094 478046 79150 478102
rect 79218 478046 79274 478102
rect 79342 478046 79398 478102
rect 78970 477922 79026 477978
rect 79094 477922 79150 477978
rect 79218 477922 79274 477978
rect 79342 477922 79398 477978
rect 78970 460294 79026 460350
rect 79094 460294 79150 460350
rect 79218 460294 79274 460350
rect 79342 460294 79398 460350
rect 78970 460170 79026 460226
rect 79094 460170 79150 460226
rect 79218 460170 79274 460226
rect 79342 460170 79398 460226
rect 78970 460046 79026 460102
rect 79094 460046 79150 460102
rect 79218 460046 79274 460102
rect 79342 460046 79398 460102
rect 78970 459922 79026 459978
rect 79094 459922 79150 459978
rect 79218 459922 79274 459978
rect 79342 459922 79398 459978
rect 78970 442294 79026 442350
rect 79094 442294 79150 442350
rect 79218 442294 79274 442350
rect 79342 442294 79398 442350
rect 78970 442170 79026 442226
rect 79094 442170 79150 442226
rect 79218 442170 79274 442226
rect 79342 442170 79398 442226
rect 78970 442046 79026 442102
rect 79094 442046 79150 442102
rect 79218 442046 79274 442102
rect 79342 442046 79398 442102
rect 78970 441922 79026 441978
rect 79094 441922 79150 441978
rect 79218 441922 79274 441978
rect 79342 441922 79398 441978
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 93250 508294 93306 508350
rect 93374 508294 93430 508350
rect 93498 508294 93554 508350
rect 93622 508294 93678 508350
rect 93250 508170 93306 508226
rect 93374 508170 93430 508226
rect 93498 508170 93554 508226
rect 93622 508170 93678 508226
rect 93250 508046 93306 508102
rect 93374 508046 93430 508102
rect 93498 508046 93554 508102
rect 93622 508046 93678 508102
rect 93250 507922 93306 507978
rect 93374 507922 93430 507978
rect 93498 507922 93554 507978
rect 93622 507922 93678 507978
rect 93250 490294 93306 490350
rect 93374 490294 93430 490350
rect 93498 490294 93554 490350
rect 93622 490294 93678 490350
rect 93250 490170 93306 490226
rect 93374 490170 93430 490226
rect 93498 490170 93554 490226
rect 93622 490170 93678 490226
rect 93250 490046 93306 490102
rect 93374 490046 93430 490102
rect 93498 490046 93554 490102
rect 93622 490046 93678 490102
rect 93250 489922 93306 489978
rect 93374 489922 93430 489978
rect 93498 489922 93554 489978
rect 93622 489922 93678 489978
rect 93250 472294 93306 472350
rect 93374 472294 93430 472350
rect 93498 472294 93554 472350
rect 93622 472294 93678 472350
rect 93250 472170 93306 472226
rect 93374 472170 93430 472226
rect 93498 472170 93554 472226
rect 93622 472170 93678 472226
rect 93250 472046 93306 472102
rect 93374 472046 93430 472102
rect 93498 472046 93554 472102
rect 93622 472046 93678 472102
rect 93250 471922 93306 471978
rect 93374 471922 93430 471978
rect 93498 471922 93554 471978
rect 93622 471922 93678 471978
rect 93250 454294 93306 454350
rect 93374 454294 93430 454350
rect 93498 454294 93554 454350
rect 93622 454294 93678 454350
rect 93250 454170 93306 454226
rect 93374 454170 93430 454226
rect 93498 454170 93554 454226
rect 93622 454170 93678 454226
rect 93250 454046 93306 454102
rect 93374 454046 93430 454102
rect 93498 454046 93554 454102
rect 93622 454046 93678 454102
rect 93250 453922 93306 453978
rect 93374 453922 93430 453978
rect 93498 453922 93554 453978
rect 93622 453922 93678 453978
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 96970 514294 97026 514350
rect 97094 514294 97150 514350
rect 97218 514294 97274 514350
rect 97342 514294 97398 514350
rect 96970 514170 97026 514226
rect 97094 514170 97150 514226
rect 97218 514170 97274 514226
rect 97342 514170 97398 514226
rect 96970 514046 97026 514102
rect 97094 514046 97150 514102
rect 97218 514046 97274 514102
rect 97342 514046 97398 514102
rect 96970 513922 97026 513978
rect 97094 513922 97150 513978
rect 97218 513922 97274 513978
rect 97342 513922 97398 513978
rect 96970 496294 97026 496350
rect 97094 496294 97150 496350
rect 97218 496294 97274 496350
rect 97342 496294 97398 496350
rect 96970 496170 97026 496226
rect 97094 496170 97150 496226
rect 97218 496170 97274 496226
rect 97342 496170 97398 496226
rect 96970 496046 97026 496102
rect 97094 496046 97150 496102
rect 97218 496046 97274 496102
rect 97342 496046 97398 496102
rect 96970 495922 97026 495978
rect 97094 495922 97150 495978
rect 97218 495922 97274 495978
rect 97342 495922 97398 495978
rect 96970 478294 97026 478350
rect 97094 478294 97150 478350
rect 97218 478294 97274 478350
rect 97342 478294 97398 478350
rect 96970 478170 97026 478226
rect 97094 478170 97150 478226
rect 97218 478170 97274 478226
rect 97342 478170 97398 478226
rect 96970 478046 97026 478102
rect 97094 478046 97150 478102
rect 97218 478046 97274 478102
rect 97342 478046 97398 478102
rect 96970 477922 97026 477978
rect 97094 477922 97150 477978
rect 97218 477922 97274 477978
rect 97342 477922 97398 477978
rect 96970 460294 97026 460350
rect 97094 460294 97150 460350
rect 97218 460294 97274 460350
rect 97342 460294 97398 460350
rect 96970 460170 97026 460226
rect 97094 460170 97150 460226
rect 97218 460170 97274 460226
rect 97342 460170 97398 460226
rect 96970 460046 97026 460102
rect 97094 460046 97150 460102
rect 97218 460046 97274 460102
rect 97342 460046 97398 460102
rect 96970 459922 97026 459978
rect 97094 459922 97150 459978
rect 97218 459922 97274 459978
rect 97342 459922 97398 459978
rect 96970 442294 97026 442350
rect 97094 442294 97150 442350
rect 97218 442294 97274 442350
rect 97342 442294 97398 442350
rect 96970 442170 97026 442226
rect 97094 442170 97150 442226
rect 97218 442170 97274 442226
rect 97342 442170 97398 442226
rect 96970 442046 97026 442102
rect 97094 442046 97150 442102
rect 97218 442046 97274 442102
rect 97342 442046 97398 442102
rect 96970 441922 97026 441978
rect 97094 441922 97150 441978
rect 97218 441922 97274 441978
rect 97342 441922 97398 441978
rect 93250 436322 93306 436378
rect 93374 436322 93430 436378
rect 93498 436322 93554 436378
rect 93622 436322 93678 436378
rect 93250 436198 93306 436254
rect 93374 436198 93430 436254
rect 93498 436198 93554 436254
rect 93622 436198 93678 436254
rect 93250 436074 93306 436130
rect 93374 436074 93430 436130
rect 93498 436074 93554 436130
rect 93622 436074 93678 436130
rect 95238 436261 95294 436317
rect 95362 436261 95418 436317
rect 95238 436137 95294 436193
rect 95362 436137 95418 436193
rect 95238 436013 95294 436069
rect 95362 436013 95418 436069
rect 64518 435889 64574 435945
rect 64642 435889 64698 435945
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 111250 508294 111306 508350
rect 111374 508294 111430 508350
rect 111498 508294 111554 508350
rect 111622 508294 111678 508350
rect 111250 508170 111306 508226
rect 111374 508170 111430 508226
rect 111498 508170 111554 508226
rect 111622 508170 111678 508226
rect 111250 508046 111306 508102
rect 111374 508046 111430 508102
rect 111498 508046 111554 508102
rect 111622 508046 111678 508102
rect 111250 507922 111306 507978
rect 111374 507922 111430 507978
rect 111498 507922 111554 507978
rect 111622 507922 111678 507978
rect 111250 490294 111306 490350
rect 111374 490294 111430 490350
rect 111498 490294 111554 490350
rect 111622 490294 111678 490350
rect 111250 490170 111306 490226
rect 111374 490170 111430 490226
rect 111498 490170 111554 490226
rect 111622 490170 111678 490226
rect 111250 490046 111306 490102
rect 111374 490046 111430 490102
rect 111498 490046 111554 490102
rect 111622 490046 111678 490102
rect 111250 489922 111306 489978
rect 111374 489922 111430 489978
rect 111498 489922 111554 489978
rect 111622 489922 111678 489978
rect 111250 472294 111306 472350
rect 111374 472294 111430 472350
rect 111498 472294 111554 472350
rect 111622 472294 111678 472350
rect 111250 472170 111306 472226
rect 111374 472170 111430 472226
rect 111498 472170 111554 472226
rect 111622 472170 111678 472226
rect 111250 472046 111306 472102
rect 111374 472046 111430 472102
rect 111498 472046 111554 472102
rect 111622 472046 111678 472102
rect 111250 471922 111306 471978
rect 111374 471922 111430 471978
rect 111498 471922 111554 471978
rect 111622 471922 111678 471978
rect 111250 454294 111306 454350
rect 111374 454294 111430 454350
rect 111498 454294 111554 454350
rect 111622 454294 111678 454350
rect 111250 454170 111306 454226
rect 111374 454170 111430 454226
rect 111498 454170 111554 454226
rect 111622 454170 111678 454226
rect 111250 454046 111306 454102
rect 111374 454046 111430 454102
rect 111498 454046 111554 454102
rect 111622 454046 111678 454102
rect 111250 453922 111306 453978
rect 111374 453922 111430 453978
rect 111498 453922 111554 453978
rect 111622 453922 111678 453978
rect 111250 436322 111306 436378
rect 111374 436322 111430 436378
rect 111498 436322 111554 436378
rect 111622 436322 111678 436378
rect 111250 436198 111306 436254
rect 111374 436198 111430 436254
rect 111498 436198 111554 436254
rect 111622 436198 111678 436254
rect 111250 436074 111306 436130
rect 111374 436074 111430 436130
rect 111498 436074 111554 436130
rect 111622 436074 111678 436130
rect 114970 598116 115026 598172
rect 115094 598116 115150 598172
rect 115218 598116 115274 598172
rect 115342 598116 115398 598172
rect 114970 597992 115026 598048
rect 115094 597992 115150 598048
rect 115218 597992 115274 598048
rect 115342 597992 115398 598048
rect 114970 597868 115026 597924
rect 115094 597868 115150 597924
rect 115218 597868 115274 597924
rect 115342 597868 115398 597924
rect 114970 597744 115026 597800
rect 115094 597744 115150 597800
rect 115218 597744 115274 597800
rect 115342 597744 115398 597800
rect 114970 586294 115026 586350
rect 115094 586294 115150 586350
rect 115218 586294 115274 586350
rect 115342 586294 115398 586350
rect 114970 586170 115026 586226
rect 115094 586170 115150 586226
rect 115218 586170 115274 586226
rect 115342 586170 115398 586226
rect 114970 586046 115026 586102
rect 115094 586046 115150 586102
rect 115218 586046 115274 586102
rect 115342 586046 115398 586102
rect 114970 585922 115026 585978
rect 115094 585922 115150 585978
rect 115218 585922 115274 585978
rect 115342 585922 115398 585978
rect 114970 568294 115026 568350
rect 115094 568294 115150 568350
rect 115218 568294 115274 568350
rect 115342 568294 115398 568350
rect 114970 568170 115026 568226
rect 115094 568170 115150 568226
rect 115218 568170 115274 568226
rect 115342 568170 115398 568226
rect 114970 568046 115026 568102
rect 115094 568046 115150 568102
rect 115218 568046 115274 568102
rect 115342 568046 115398 568102
rect 114970 567922 115026 567978
rect 115094 567922 115150 567978
rect 115218 567922 115274 567978
rect 115342 567922 115398 567978
rect 114970 550294 115026 550350
rect 115094 550294 115150 550350
rect 115218 550294 115274 550350
rect 115342 550294 115398 550350
rect 114970 550170 115026 550226
rect 115094 550170 115150 550226
rect 115218 550170 115274 550226
rect 115342 550170 115398 550226
rect 114970 550046 115026 550102
rect 115094 550046 115150 550102
rect 115218 550046 115274 550102
rect 115342 550046 115398 550102
rect 114970 549922 115026 549978
rect 115094 549922 115150 549978
rect 115218 549922 115274 549978
rect 115342 549922 115398 549978
rect 114970 532294 115026 532350
rect 115094 532294 115150 532350
rect 115218 532294 115274 532350
rect 115342 532294 115398 532350
rect 114970 532170 115026 532226
rect 115094 532170 115150 532226
rect 115218 532170 115274 532226
rect 115342 532170 115398 532226
rect 114970 532046 115026 532102
rect 115094 532046 115150 532102
rect 115218 532046 115274 532102
rect 115342 532046 115398 532102
rect 114970 531922 115026 531978
rect 115094 531922 115150 531978
rect 115218 531922 115274 531978
rect 115342 531922 115398 531978
rect 114970 514294 115026 514350
rect 115094 514294 115150 514350
rect 115218 514294 115274 514350
rect 115342 514294 115398 514350
rect 114970 514170 115026 514226
rect 115094 514170 115150 514226
rect 115218 514170 115274 514226
rect 115342 514170 115398 514226
rect 114970 514046 115026 514102
rect 115094 514046 115150 514102
rect 115218 514046 115274 514102
rect 115342 514046 115398 514102
rect 114970 513922 115026 513978
rect 115094 513922 115150 513978
rect 115218 513922 115274 513978
rect 115342 513922 115398 513978
rect 114970 496294 115026 496350
rect 115094 496294 115150 496350
rect 115218 496294 115274 496350
rect 115342 496294 115398 496350
rect 114970 496170 115026 496226
rect 115094 496170 115150 496226
rect 115218 496170 115274 496226
rect 115342 496170 115398 496226
rect 114970 496046 115026 496102
rect 115094 496046 115150 496102
rect 115218 496046 115274 496102
rect 115342 496046 115398 496102
rect 114970 495922 115026 495978
rect 115094 495922 115150 495978
rect 115218 495922 115274 495978
rect 115342 495922 115398 495978
rect 114970 478294 115026 478350
rect 115094 478294 115150 478350
rect 115218 478294 115274 478350
rect 115342 478294 115398 478350
rect 114970 478170 115026 478226
rect 115094 478170 115150 478226
rect 115218 478170 115274 478226
rect 115342 478170 115398 478226
rect 114970 478046 115026 478102
rect 115094 478046 115150 478102
rect 115218 478046 115274 478102
rect 115342 478046 115398 478102
rect 114970 477922 115026 477978
rect 115094 477922 115150 477978
rect 115218 477922 115274 477978
rect 115342 477922 115398 477978
rect 114970 460294 115026 460350
rect 115094 460294 115150 460350
rect 115218 460294 115274 460350
rect 115342 460294 115398 460350
rect 114970 460170 115026 460226
rect 115094 460170 115150 460226
rect 115218 460170 115274 460226
rect 115342 460170 115398 460226
rect 114970 460046 115026 460102
rect 115094 460046 115150 460102
rect 115218 460046 115274 460102
rect 115342 460046 115398 460102
rect 114970 459922 115026 459978
rect 115094 459922 115150 459978
rect 115218 459922 115274 459978
rect 115342 459922 115398 459978
rect 114970 442294 115026 442350
rect 115094 442294 115150 442350
rect 115218 442294 115274 442350
rect 115342 442294 115398 442350
rect 114970 442170 115026 442226
rect 115094 442170 115150 442226
rect 115218 442170 115274 442226
rect 115342 442170 115398 442226
rect 114970 442046 115026 442102
rect 115094 442046 115150 442102
rect 115218 442046 115274 442102
rect 115342 442046 115398 442102
rect 114970 441922 115026 441978
rect 115094 441922 115150 441978
rect 115218 441922 115274 441978
rect 115342 441922 115398 441978
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 129250 526294 129306 526350
rect 129374 526294 129430 526350
rect 129498 526294 129554 526350
rect 129622 526294 129678 526350
rect 129250 526170 129306 526226
rect 129374 526170 129430 526226
rect 129498 526170 129554 526226
rect 129622 526170 129678 526226
rect 129250 526046 129306 526102
rect 129374 526046 129430 526102
rect 129498 526046 129554 526102
rect 129622 526046 129678 526102
rect 129250 525922 129306 525978
rect 129374 525922 129430 525978
rect 129498 525922 129554 525978
rect 129622 525922 129678 525978
rect 129250 508294 129306 508350
rect 129374 508294 129430 508350
rect 129498 508294 129554 508350
rect 129622 508294 129678 508350
rect 129250 508170 129306 508226
rect 129374 508170 129430 508226
rect 129498 508170 129554 508226
rect 129622 508170 129678 508226
rect 129250 508046 129306 508102
rect 129374 508046 129430 508102
rect 129498 508046 129554 508102
rect 129622 508046 129678 508102
rect 129250 507922 129306 507978
rect 129374 507922 129430 507978
rect 129498 507922 129554 507978
rect 129622 507922 129678 507978
rect 129250 490294 129306 490350
rect 129374 490294 129430 490350
rect 129498 490294 129554 490350
rect 129622 490294 129678 490350
rect 129250 490170 129306 490226
rect 129374 490170 129430 490226
rect 129498 490170 129554 490226
rect 129622 490170 129678 490226
rect 129250 490046 129306 490102
rect 129374 490046 129430 490102
rect 129498 490046 129554 490102
rect 129622 490046 129678 490102
rect 129250 489922 129306 489978
rect 129374 489922 129430 489978
rect 129498 489922 129554 489978
rect 129622 489922 129678 489978
rect 129250 472294 129306 472350
rect 129374 472294 129430 472350
rect 129498 472294 129554 472350
rect 129622 472294 129678 472350
rect 129250 472170 129306 472226
rect 129374 472170 129430 472226
rect 129498 472170 129554 472226
rect 129622 472170 129678 472226
rect 129250 472046 129306 472102
rect 129374 472046 129430 472102
rect 129498 472046 129554 472102
rect 129622 472046 129678 472102
rect 129250 471922 129306 471978
rect 129374 471922 129430 471978
rect 129498 471922 129554 471978
rect 129622 471922 129678 471978
rect 129250 454294 129306 454350
rect 129374 454294 129430 454350
rect 129498 454294 129554 454350
rect 129622 454294 129678 454350
rect 129250 454170 129306 454226
rect 129374 454170 129430 454226
rect 129498 454170 129554 454226
rect 129622 454170 129678 454226
rect 129250 454046 129306 454102
rect 129374 454046 129430 454102
rect 129498 454046 129554 454102
rect 129622 454046 129678 454102
rect 129250 453922 129306 453978
rect 129374 453922 129430 453978
rect 129498 453922 129554 453978
rect 129622 453922 129678 453978
rect 125958 436261 126014 436317
rect 126082 436261 126138 436317
rect 125958 436137 126014 436193
rect 126082 436137 126138 436193
rect 125958 436013 126014 436069
rect 126082 436013 126138 436069
rect 95238 435889 95294 435945
rect 95362 435889 95418 435945
rect 129250 436322 129306 436378
rect 129374 436322 129430 436378
rect 129498 436322 129554 436378
rect 129622 436322 129678 436378
rect 129250 436198 129306 436254
rect 129374 436198 129430 436254
rect 129498 436198 129554 436254
rect 129622 436198 129678 436254
rect 129250 436074 129306 436130
rect 129374 436074 129430 436130
rect 129498 436074 129554 436130
rect 129622 436074 129678 436130
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 132970 514294 133026 514350
rect 133094 514294 133150 514350
rect 133218 514294 133274 514350
rect 133342 514294 133398 514350
rect 132970 514170 133026 514226
rect 133094 514170 133150 514226
rect 133218 514170 133274 514226
rect 133342 514170 133398 514226
rect 132970 514046 133026 514102
rect 133094 514046 133150 514102
rect 133218 514046 133274 514102
rect 133342 514046 133398 514102
rect 132970 513922 133026 513978
rect 133094 513922 133150 513978
rect 133218 513922 133274 513978
rect 133342 513922 133398 513978
rect 132970 496294 133026 496350
rect 133094 496294 133150 496350
rect 133218 496294 133274 496350
rect 133342 496294 133398 496350
rect 132970 496170 133026 496226
rect 133094 496170 133150 496226
rect 133218 496170 133274 496226
rect 133342 496170 133398 496226
rect 132970 496046 133026 496102
rect 133094 496046 133150 496102
rect 133218 496046 133274 496102
rect 133342 496046 133398 496102
rect 132970 495922 133026 495978
rect 133094 495922 133150 495978
rect 133218 495922 133274 495978
rect 133342 495922 133398 495978
rect 132970 478294 133026 478350
rect 133094 478294 133150 478350
rect 133218 478294 133274 478350
rect 133342 478294 133398 478350
rect 132970 478170 133026 478226
rect 133094 478170 133150 478226
rect 133218 478170 133274 478226
rect 133342 478170 133398 478226
rect 132970 478046 133026 478102
rect 133094 478046 133150 478102
rect 133218 478046 133274 478102
rect 133342 478046 133398 478102
rect 132970 477922 133026 477978
rect 133094 477922 133150 477978
rect 133218 477922 133274 477978
rect 133342 477922 133398 477978
rect 132970 460294 133026 460350
rect 133094 460294 133150 460350
rect 133218 460294 133274 460350
rect 133342 460294 133398 460350
rect 132970 460170 133026 460226
rect 133094 460170 133150 460226
rect 133218 460170 133274 460226
rect 133342 460170 133398 460226
rect 132970 460046 133026 460102
rect 133094 460046 133150 460102
rect 133218 460046 133274 460102
rect 133342 460046 133398 460102
rect 132970 459922 133026 459978
rect 133094 459922 133150 459978
rect 133218 459922 133274 459978
rect 133342 459922 133398 459978
rect 132970 442294 133026 442350
rect 133094 442294 133150 442350
rect 133218 442294 133274 442350
rect 133342 442294 133398 442350
rect 132970 442170 133026 442226
rect 133094 442170 133150 442226
rect 133218 442170 133274 442226
rect 133342 442170 133398 442226
rect 132970 442046 133026 442102
rect 133094 442046 133150 442102
rect 133218 442046 133274 442102
rect 133342 442046 133398 442102
rect 132970 441922 133026 441978
rect 133094 441922 133150 441978
rect 133218 441922 133274 441978
rect 133342 441922 133398 441978
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 147250 526294 147306 526350
rect 147374 526294 147430 526350
rect 147498 526294 147554 526350
rect 147622 526294 147678 526350
rect 147250 526170 147306 526226
rect 147374 526170 147430 526226
rect 147498 526170 147554 526226
rect 147622 526170 147678 526226
rect 147250 526046 147306 526102
rect 147374 526046 147430 526102
rect 147498 526046 147554 526102
rect 147622 526046 147678 526102
rect 147250 525922 147306 525978
rect 147374 525922 147430 525978
rect 147498 525922 147554 525978
rect 147622 525922 147678 525978
rect 147250 508294 147306 508350
rect 147374 508294 147430 508350
rect 147498 508294 147554 508350
rect 147622 508294 147678 508350
rect 147250 508170 147306 508226
rect 147374 508170 147430 508226
rect 147498 508170 147554 508226
rect 147622 508170 147678 508226
rect 147250 508046 147306 508102
rect 147374 508046 147430 508102
rect 147498 508046 147554 508102
rect 147622 508046 147678 508102
rect 147250 507922 147306 507978
rect 147374 507922 147430 507978
rect 147498 507922 147554 507978
rect 147622 507922 147678 507978
rect 147250 490294 147306 490350
rect 147374 490294 147430 490350
rect 147498 490294 147554 490350
rect 147622 490294 147678 490350
rect 147250 490170 147306 490226
rect 147374 490170 147430 490226
rect 147498 490170 147554 490226
rect 147622 490170 147678 490226
rect 147250 490046 147306 490102
rect 147374 490046 147430 490102
rect 147498 490046 147554 490102
rect 147622 490046 147678 490102
rect 147250 489922 147306 489978
rect 147374 489922 147430 489978
rect 147498 489922 147554 489978
rect 147622 489922 147678 489978
rect 147250 472294 147306 472350
rect 147374 472294 147430 472350
rect 147498 472294 147554 472350
rect 147622 472294 147678 472350
rect 147250 472170 147306 472226
rect 147374 472170 147430 472226
rect 147498 472170 147554 472226
rect 147622 472170 147678 472226
rect 147250 472046 147306 472102
rect 147374 472046 147430 472102
rect 147498 472046 147554 472102
rect 147622 472046 147678 472102
rect 147250 471922 147306 471978
rect 147374 471922 147430 471978
rect 147498 471922 147554 471978
rect 147622 471922 147678 471978
rect 147250 454294 147306 454350
rect 147374 454294 147430 454350
rect 147498 454294 147554 454350
rect 147622 454294 147678 454350
rect 147250 454170 147306 454226
rect 147374 454170 147430 454226
rect 147498 454170 147554 454226
rect 147622 454170 147678 454226
rect 147250 454046 147306 454102
rect 147374 454046 147430 454102
rect 147498 454046 147554 454102
rect 147622 454046 147678 454102
rect 147250 453922 147306 453978
rect 147374 453922 147430 453978
rect 147498 453922 147554 453978
rect 147622 453922 147678 453978
rect 147250 436322 147306 436378
rect 147374 436322 147430 436378
rect 147498 436322 147554 436378
rect 147622 436322 147678 436378
rect 147250 436198 147306 436254
rect 147374 436198 147430 436254
rect 147498 436198 147554 436254
rect 147622 436198 147678 436254
rect 147250 436074 147306 436130
rect 147374 436074 147430 436130
rect 147498 436074 147554 436130
rect 147622 436074 147678 436130
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 150970 514294 151026 514350
rect 151094 514294 151150 514350
rect 151218 514294 151274 514350
rect 151342 514294 151398 514350
rect 150970 514170 151026 514226
rect 151094 514170 151150 514226
rect 151218 514170 151274 514226
rect 151342 514170 151398 514226
rect 150970 514046 151026 514102
rect 151094 514046 151150 514102
rect 151218 514046 151274 514102
rect 151342 514046 151398 514102
rect 150970 513922 151026 513978
rect 151094 513922 151150 513978
rect 151218 513922 151274 513978
rect 151342 513922 151398 513978
rect 150970 496294 151026 496350
rect 151094 496294 151150 496350
rect 151218 496294 151274 496350
rect 151342 496294 151398 496350
rect 150970 496170 151026 496226
rect 151094 496170 151150 496226
rect 151218 496170 151274 496226
rect 151342 496170 151398 496226
rect 150970 496046 151026 496102
rect 151094 496046 151150 496102
rect 151218 496046 151274 496102
rect 151342 496046 151398 496102
rect 150970 495922 151026 495978
rect 151094 495922 151150 495978
rect 151218 495922 151274 495978
rect 151342 495922 151398 495978
rect 150970 478294 151026 478350
rect 151094 478294 151150 478350
rect 151218 478294 151274 478350
rect 151342 478294 151398 478350
rect 150970 478170 151026 478226
rect 151094 478170 151150 478226
rect 151218 478170 151274 478226
rect 151342 478170 151398 478226
rect 150970 478046 151026 478102
rect 151094 478046 151150 478102
rect 151218 478046 151274 478102
rect 151342 478046 151398 478102
rect 150970 477922 151026 477978
rect 151094 477922 151150 477978
rect 151218 477922 151274 477978
rect 151342 477922 151398 477978
rect 150970 460294 151026 460350
rect 151094 460294 151150 460350
rect 151218 460294 151274 460350
rect 151342 460294 151398 460350
rect 150970 460170 151026 460226
rect 151094 460170 151150 460226
rect 151218 460170 151274 460226
rect 151342 460170 151398 460226
rect 150970 460046 151026 460102
rect 151094 460046 151150 460102
rect 151218 460046 151274 460102
rect 151342 460046 151398 460102
rect 150970 459922 151026 459978
rect 151094 459922 151150 459978
rect 151218 459922 151274 459978
rect 151342 459922 151398 459978
rect 150970 442294 151026 442350
rect 151094 442294 151150 442350
rect 151218 442294 151274 442350
rect 151342 442294 151398 442350
rect 150970 442170 151026 442226
rect 151094 442170 151150 442226
rect 151218 442170 151274 442226
rect 151342 442170 151398 442226
rect 150970 442046 151026 442102
rect 151094 442046 151150 442102
rect 151218 442046 151274 442102
rect 151342 442046 151398 442102
rect 150970 441922 151026 441978
rect 151094 441922 151150 441978
rect 151218 441922 151274 441978
rect 151342 441922 151398 441978
rect 165250 597156 165306 597212
rect 165374 597156 165430 597212
rect 165498 597156 165554 597212
rect 165622 597156 165678 597212
rect 165250 597032 165306 597088
rect 165374 597032 165430 597088
rect 165498 597032 165554 597088
rect 165622 597032 165678 597088
rect 165250 596908 165306 596964
rect 165374 596908 165430 596964
rect 165498 596908 165554 596964
rect 165622 596908 165678 596964
rect 165250 596784 165306 596840
rect 165374 596784 165430 596840
rect 165498 596784 165554 596840
rect 165622 596784 165678 596840
rect 165250 580294 165306 580350
rect 165374 580294 165430 580350
rect 165498 580294 165554 580350
rect 165622 580294 165678 580350
rect 165250 580170 165306 580226
rect 165374 580170 165430 580226
rect 165498 580170 165554 580226
rect 165622 580170 165678 580226
rect 165250 580046 165306 580102
rect 165374 580046 165430 580102
rect 165498 580046 165554 580102
rect 165622 580046 165678 580102
rect 165250 579922 165306 579978
rect 165374 579922 165430 579978
rect 165498 579922 165554 579978
rect 165622 579922 165678 579978
rect 165250 562294 165306 562350
rect 165374 562294 165430 562350
rect 165498 562294 165554 562350
rect 165622 562294 165678 562350
rect 165250 562170 165306 562226
rect 165374 562170 165430 562226
rect 165498 562170 165554 562226
rect 165622 562170 165678 562226
rect 165250 562046 165306 562102
rect 165374 562046 165430 562102
rect 165498 562046 165554 562102
rect 165622 562046 165678 562102
rect 165250 561922 165306 561978
rect 165374 561922 165430 561978
rect 165498 561922 165554 561978
rect 165622 561922 165678 561978
rect 165250 544294 165306 544350
rect 165374 544294 165430 544350
rect 165498 544294 165554 544350
rect 165622 544294 165678 544350
rect 165250 544170 165306 544226
rect 165374 544170 165430 544226
rect 165498 544170 165554 544226
rect 165622 544170 165678 544226
rect 165250 544046 165306 544102
rect 165374 544046 165430 544102
rect 165498 544046 165554 544102
rect 165622 544046 165678 544102
rect 165250 543922 165306 543978
rect 165374 543922 165430 543978
rect 165498 543922 165554 543978
rect 165622 543922 165678 543978
rect 165250 526294 165306 526350
rect 165374 526294 165430 526350
rect 165498 526294 165554 526350
rect 165622 526294 165678 526350
rect 165250 526170 165306 526226
rect 165374 526170 165430 526226
rect 165498 526170 165554 526226
rect 165622 526170 165678 526226
rect 165250 526046 165306 526102
rect 165374 526046 165430 526102
rect 165498 526046 165554 526102
rect 165622 526046 165678 526102
rect 165250 525922 165306 525978
rect 165374 525922 165430 525978
rect 165498 525922 165554 525978
rect 165622 525922 165678 525978
rect 165250 508294 165306 508350
rect 165374 508294 165430 508350
rect 165498 508294 165554 508350
rect 165622 508294 165678 508350
rect 165250 508170 165306 508226
rect 165374 508170 165430 508226
rect 165498 508170 165554 508226
rect 165622 508170 165678 508226
rect 165250 508046 165306 508102
rect 165374 508046 165430 508102
rect 165498 508046 165554 508102
rect 165622 508046 165678 508102
rect 165250 507922 165306 507978
rect 165374 507922 165430 507978
rect 165498 507922 165554 507978
rect 165622 507922 165678 507978
rect 165250 490294 165306 490350
rect 165374 490294 165430 490350
rect 165498 490294 165554 490350
rect 165622 490294 165678 490350
rect 165250 490170 165306 490226
rect 165374 490170 165430 490226
rect 165498 490170 165554 490226
rect 165622 490170 165678 490226
rect 165250 490046 165306 490102
rect 165374 490046 165430 490102
rect 165498 490046 165554 490102
rect 165622 490046 165678 490102
rect 165250 489922 165306 489978
rect 165374 489922 165430 489978
rect 165498 489922 165554 489978
rect 165622 489922 165678 489978
rect 165250 472294 165306 472350
rect 165374 472294 165430 472350
rect 165498 472294 165554 472350
rect 165622 472294 165678 472350
rect 165250 472170 165306 472226
rect 165374 472170 165430 472226
rect 165498 472170 165554 472226
rect 165622 472170 165678 472226
rect 165250 472046 165306 472102
rect 165374 472046 165430 472102
rect 165498 472046 165554 472102
rect 165622 472046 165678 472102
rect 165250 471922 165306 471978
rect 165374 471922 165430 471978
rect 165498 471922 165554 471978
rect 165622 471922 165678 471978
rect 165250 454294 165306 454350
rect 165374 454294 165430 454350
rect 165498 454294 165554 454350
rect 165622 454294 165678 454350
rect 165250 454170 165306 454226
rect 165374 454170 165430 454226
rect 165498 454170 165554 454226
rect 165622 454170 165678 454226
rect 165250 454046 165306 454102
rect 165374 454046 165430 454102
rect 165498 454046 165554 454102
rect 165622 454046 165678 454102
rect 165250 453922 165306 453978
rect 165374 453922 165430 453978
rect 165498 453922 165554 453978
rect 165622 453922 165678 453978
rect 156678 436261 156734 436317
rect 156802 436261 156858 436317
rect 156678 436137 156734 436193
rect 156802 436137 156858 436193
rect 156678 436013 156734 436069
rect 156802 436013 156858 436069
rect 125958 435889 126014 435945
rect 126082 435889 126138 435945
rect 165250 436322 165306 436378
rect 165374 436322 165430 436378
rect 165498 436322 165554 436378
rect 165622 436322 165678 436378
rect 165250 436198 165306 436254
rect 165374 436198 165430 436254
rect 165498 436198 165554 436254
rect 165622 436198 165678 436254
rect 165250 436074 165306 436130
rect 165374 436074 165430 436130
rect 165498 436074 165554 436130
rect 165622 436074 165678 436130
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 168970 514294 169026 514350
rect 169094 514294 169150 514350
rect 169218 514294 169274 514350
rect 169342 514294 169398 514350
rect 168970 514170 169026 514226
rect 169094 514170 169150 514226
rect 169218 514170 169274 514226
rect 169342 514170 169398 514226
rect 168970 514046 169026 514102
rect 169094 514046 169150 514102
rect 169218 514046 169274 514102
rect 169342 514046 169398 514102
rect 168970 513922 169026 513978
rect 169094 513922 169150 513978
rect 169218 513922 169274 513978
rect 169342 513922 169398 513978
rect 168970 496294 169026 496350
rect 169094 496294 169150 496350
rect 169218 496294 169274 496350
rect 169342 496294 169398 496350
rect 168970 496170 169026 496226
rect 169094 496170 169150 496226
rect 169218 496170 169274 496226
rect 169342 496170 169398 496226
rect 168970 496046 169026 496102
rect 169094 496046 169150 496102
rect 169218 496046 169274 496102
rect 169342 496046 169398 496102
rect 168970 495922 169026 495978
rect 169094 495922 169150 495978
rect 169218 495922 169274 495978
rect 169342 495922 169398 495978
rect 168970 478294 169026 478350
rect 169094 478294 169150 478350
rect 169218 478294 169274 478350
rect 169342 478294 169398 478350
rect 168970 478170 169026 478226
rect 169094 478170 169150 478226
rect 169218 478170 169274 478226
rect 169342 478170 169398 478226
rect 168970 478046 169026 478102
rect 169094 478046 169150 478102
rect 169218 478046 169274 478102
rect 169342 478046 169398 478102
rect 168970 477922 169026 477978
rect 169094 477922 169150 477978
rect 169218 477922 169274 477978
rect 169342 477922 169398 477978
rect 168970 460294 169026 460350
rect 169094 460294 169150 460350
rect 169218 460294 169274 460350
rect 169342 460294 169398 460350
rect 168970 460170 169026 460226
rect 169094 460170 169150 460226
rect 169218 460170 169274 460226
rect 169342 460170 169398 460226
rect 168970 460046 169026 460102
rect 169094 460046 169150 460102
rect 169218 460046 169274 460102
rect 169342 460046 169398 460102
rect 168970 459922 169026 459978
rect 169094 459922 169150 459978
rect 169218 459922 169274 459978
rect 169342 459922 169398 459978
rect 168970 442294 169026 442350
rect 169094 442294 169150 442350
rect 169218 442294 169274 442350
rect 169342 442294 169398 442350
rect 168970 442170 169026 442226
rect 169094 442170 169150 442226
rect 169218 442170 169274 442226
rect 169342 442170 169398 442226
rect 168970 442046 169026 442102
rect 169094 442046 169150 442102
rect 169218 442046 169274 442102
rect 169342 442046 169398 442102
rect 168970 441922 169026 441978
rect 169094 441922 169150 441978
rect 169218 441922 169274 441978
rect 169342 441922 169398 441978
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 183250 526294 183306 526350
rect 183374 526294 183430 526350
rect 183498 526294 183554 526350
rect 183622 526294 183678 526350
rect 183250 526170 183306 526226
rect 183374 526170 183430 526226
rect 183498 526170 183554 526226
rect 183622 526170 183678 526226
rect 183250 526046 183306 526102
rect 183374 526046 183430 526102
rect 183498 526046 183554 526102
rect 183622 526046 183678 526102
rect 183250 525922 183306 525978
rect 183374 525922 183430 525978
rect 183498 525922 183554 525978
rect 183622 525922 183678 525978
rect 183250 508294 183306 508350
rect 183374 508294 183430 508350
rect 183498 508294 183554 508350
rect 183622 508294 183678 508350
rect 183250 508170 183306 508226
rect 183374 508170 183430 508226
rect 183498 508170 183554 508226
rect 183622 508170 183678 508226
rect 183250 508046 183306 508102
rect 183374 508046 183430 508102
rect 183498 508046 183554 508102
rect 183622 508046 183678 508102
rect 183250 507922 183306 507978
rect 183374 507922 183430 507978
rect 183498 507922 183554 507978
rect 183622 507922 183678 507978
rect 183250 490294 183306 490350
rect 183374 490294 183430 490350
rect 183498 490294 183554 490350
rect 183622 490294 183678 490350
rect 183250 490170 183306 490226
rect 183374 490170 183430 490226
rect 183498 490170 183554 490226
rect 183622 490170 183678 490226
rect 183250 490046 183306 490102
rect 183374 490046 183430 490102
rect 183498 490046 183554 490102
rect 183622 490046 183678 490102
rect 183250 489922 183306 489978
rect 183374 489922 183430 489978
rect 183498 489922 183554 489978
rect 183622 489922 183678 489978
rect 183250 472294 183306 472350
rect 183374 472294 183430 472350
rect 183498 472294 183554 472350
rect 183622 472294 183678 472350
rect 183250 472170 183306 472226
rect 183374 472170 183430 472226
rect 183498 472170 183554 472226
rect 183622 472170 183678 472226
rect 183250 472046 183306 472102
rect 183374 472046 183430 472102
rect 183498 472046 183554 472102
rect 183622 472046 183678 472102
rect 183250 471922 183306 471978
rect 183374 471922 183430 471978
rect 183498 471922 183554 471978
rect 183622 471922 183678 471978
rect 183250 454294 183306 454350
rect 183374 454294 183430 454350
rect 183498 454294 183554 454350
rect 183622 454294 183678 454350
rect 183250 454170 183306 454226
rect 183374 454170 183430 454226
rect 183498 454170 183554 454226
rect 183622 454170 183678 454226
rect 183250 454046 183306 454102
rect 183374 454046 183430 454102
rect 183498 454046 183554 454102
rect 183622 454046 183678 454102
rect 183250 453922 183306 453978
rect 183374 453922 183430 453978
rect 183498 453922 183554 453978
rect 183622 453922 183678 453978
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 186970 514294 187026 514350
rect 187094 514294 187150 514350
rect 187218 514294 187274 514350
rect 187342 514294 187398 514350
rect 186970 514170 187026 514226
rect 187094 514170 187150 514226
rect 187218 514170 187274 514226
rect 187342 514170 187398 514226
rect 186970 514046 187026 514102
rect 187094 514046 187150 514102
rect 187218 514046 187274 514102
rect 187342 514046 187398 514102
rect 186970 513922 187026 513978
rect 187094 513922 187150 513978
rect 187218 513922 187274 513978
rect 187342 513922 187398 513978
rect 186970 496294 187026 496350
rect 187094 496294 187150 496350
rect 187218 496294 187274 496350
rect 187342 496294 187398 496350
rect 186970 496170 187026 496226
rect 187094 496170 187150 496226
rect 187218 496170 187274 496226
rect 187342 496170 187398 496226
rect 186970 496046 187026 496102
rect 187094 496046 187150 496102
rect 187218 496046 187274 496102
rect 187342 496046 187398 496102
rect 186970 495922 187026 495978
rect 187094 495922 187150 495978
rect 187218 495922 187274 495978
rect 187342 495922 187398 495978
rect 186970 478294 187026 478350
rect 187094 478294 187150 478350
rect 187218 478294 187274 478350
rect 187342 478294 187398 478350
rect 186970 478170 187026 478226
rect 187094 478170 187150 478226
rect 187218 478170 187274 478226
rect 187342 478170 187398 478226
rect 186970 478046 187026 478102
rect 187094 478046 187150 478102
rect 187218 478046 187274 478102
rect 187342 478046 187398 478102
rect 186970 477922 187026 477978
rect 187094 477922 187150 477978
rect 187218 477922 187274 477978
rect 187342 477922 187398 477978
rect 186970 460294 187026 460350
rect 187094 460294 187150 460350
rect 187218 460294 187274 460350
rect 187342 460294 187398 460350
rect 186970 460170 187026 460226
rect 187094 460170 187150 460226
rect 187218 460170 187274 460226
rect 187342 460170 187398 460226
rect 186970 460046 187026 460102
rect 187094 460046 187150 460102
rect 187218 460046 187274 460102
rect 187342 460046 187398 460102
rect 186970 459922 187026 459978
rect 187094 459922 187150 459978
rect 187218 459922 187274 459978
rect 187342 459922 187398 459978
rect 186970 442294 187026 442350
rect 187094 442294 187150 442350
rect 187218 442294 187274 442350
rect 187342 442294 187398 442350
rect 186970 442170 187026 442226
rect 187094 442170 187150 442226
rect 187218 442170 187274 442226
rect 187342 442170 187398 442226
rect 186970 442046 187026 442102
rect 187094 442046 187150 442102
rect 187218 442046 187274 442102
rect 187342 442046 187398 442102
rect 186970 441922 187026 441978
rect 187094 441922 187150 441978
rect 187218 441922 187274 441978
rect 187342 441922 187398 441978
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 201250 526294 201306 526350
rect 201374 526294 201430 526350
rect 201498 526294 201554 526350
rect 201622 526294 201678 526350
rect 201250 526170 201306 526226
rect 201374 526170 201430 526226
rect 201498 526170 201554 526226
rect 201622 526170 201678 526226
rect 201250 526046 201306 526102
rect 201374 526046 201430 526102
rect 201498 526046 201554 526102
rect 201622 526046 201678 526102
rect 201250 525922 201306 525978
rect 201374 525922 201430 525978
rect 201498 525922 201554 525978
rect 201622 525922 201678 525978
rect 201250 508294 201306 508350
rect 201374 508294 201430 508350
rect 201498 508294 201554 508350
rect 201622 508294 201678 508350
rect 201250 508170 201306 508226
rect 201374 508170 201430 508226
rect 201498 508170 201554 508226
rect 201622 508170 201678 508226
rect 201250 508046 201306 508102
rect 201374 508046 201430 508102
rect 201498 508046 201554 508102
rect 201622 508046 201678 508102
rect 201250 507922 201306 507978
rect 201374 507922 201430 507978
rect 201498 507922 201554 507978
rect 201622 507922 201678 507978
rect 201250 490294 201306 490350
rect 201374 490294 201430 490350
rect 201498 490294 201554 490350
rect 201622 490294 201678 490350
rect 201250 490170 201306 490226
rect 201374 490170 201430 490226
rect 201498 490170 201554 490226
rect 201622 490170 201678 490226
rect 201250 490046 201306 490102
rect 201374 490046 201430 490102
rect 201498 490046 201554 490102
rect 201622 490046 201678 490102
rect 201250 489922 201306 489978
rect 201374 489922 201430 489978
rect 201498 489922 201554 489978
rect 201622 489922 201678 489978
rect 201250 472294 201306 472350
rect 201374 472294 201430 472350
rect 201498 472294 201554 472350
rect 201622 472294 201678 472350
rect 201250 472170 201306 472226
rect 201374 472170 201430 472226
rect 201498 472170 201554 472226
rect 201622 472170 201678 472226
rect 201250 472046 201306 472102
rect 201374 472046 201430 472102
rect 201498 472046 201554 472102
rect 201622 472046 201678 472102
rect 201250 471922 201306 471978
rect 201374 471922 201430 471978
rect 201498 471922 201554 471978
rect 201622 471922 201678 471978
rect 201250 454294 201306 454350
rect 201374 454294 201430 454350
rect 201498 454294 201554 454350
rect 201622 454294 201678 454350
rect 201250 454170 201306 454226
rect 201374 454170 201430 454226
rect 201498 454170 201554 454226
rect 201622 454170 201678 454226
rect 201250 454046 201306 454102
rect 201374 454046 201430 454102
rect 201498 454046 201554 454102
rect 201622 454046 201678 454102
rect 201250 453922 201306 453978
rect 201374 453922 201430 453978
rect 201498 453922 201554 453978
rect 201622 453922 201678 453978
rect 183250 436322 183306 436378
rect 183374 436322 183430 436378
rect 183498 436322 183554 436378
rect 183622 436322 183678 436378
rect 183250 436198 183306 436254
rect 183374 436198 183430 436254
rect 183498 436198 183554 436254
rect 183622 436198 183678 436254
rect 183250 436074 183306 436130
rect 183374 436074 183430 436130
rect 183498 436074 183554 436130
rect 183622 436074 183678 436130
rect 187398 436261 187454 436317
rect 187522 436261 187578 436317
rect 187398 436137 187454 436193
rect 187522 436137 187578 436193
rect 187398 436013 187454 436069
rect 187522 436013 187578 436069
rect 156678 435889 156734 435945
rect 156802 435889 156858 435945
rect 201250 436322 201306 436378
rect 201374 436322 201430 436378
rect 201498 436322 201554 436378
rect 201622 436322 201678 436378
rect 201250 436198 201306 436254
rect 201374 436198 201430 436254
rect 201498 436198 201554 436254
rect 201622 436198 201678 436254
rect 201250 436074 201306 436130
rect 201374 436074 201430 436130
rect 201498 436074 201554 436130
rect 201622 436074 201678 436130
rect 204970 598116 205026 598172
rect 205094 598116 205150 598172
rect 205218 598116 205274 598172
rect 205342 598116 205398 598172
rect 204970 597992 205026 598048
rect 205094 597992 205150 598048
rect 205218 597992 205274 598048
rect 205342 597992 205398 598048
rect 204970 597868 205026 597924
rect 205094 597868 205150 597924
rect 205218 597868 205274 597924
rect 205342 597868 205398 597924
rect 204970 597744 205026 597800
rect 205094 597744 205150 597800
rect 205218 597744 205274 597800
rect 205342 597744 205398 597800
rect 204970 586294 205026 586350
rect 205094 586294 205150 586350
rect 205218 586294 205274 586350
rect 205342 586294 205398 586350
rect 204970 586170 205026 586226
rect 205094 586170 205150 586226
rect 205218 586170 205274 586226
rect 205342 586170 205398 586226
rect 204970 586046 205026 586102
rect 205094 586046 205150 586102
rect 205218 586046 205274 586102
rect 205342 586046 205398 586102
rect 204970 585922 205026 585978
rect 205094 585922 205150 585978
rect 205218 585922 205274 585978
rect 205342 585922 205398 585978
rect 204970 568294 205026 568350
rect 205094 568294 205150 568350
rect 205218 568294 205274 568350
rect 205342 568294 205398 568350
rect 204970 568170 205026 568226
rect 205094 568170 205150 568226
rect 205218 568170 205274 568226
rect 205342 568170 205398 568226
rect 204970 568046 205026 568102
rect 205094 568046 205150 568102
rect 205218 568046 205274 568102
rect 205342 568046 205398 568102
rect 204970 567922 205026 567978
rect 205094 567922 205150 567978
rect 205218 567922 205274 567978
rect 205342 567922 205398 567978
rect 204970 550294 205026 550350
rect 205094 550294 205150 550350
rect 205218 550294 205274 550350
rect 205342 550294 205398 550350
rect 204970 550170 205026 550226
rect 205094 550170 205150 550226
rect 205218 550170 205274 550226
rect 205342 550170 205398 550226
rect 204970 550046 205026 550102
rect 205094 550046 205150 550102
rect 205218 550046 205274 550102
rect 205342 550046 205398 550102
rect 204970 549922 205026 549978
rect 205094 549922 205150 549978
rect 205218 549922 205274 549978
rect 205342 549922 205398 549978
rect 204970 532294 205026 532350
rect 205094 532294 205150 532350
rect 205218 532294 205274 532350
rect 205342 532294 205398 532350
rect 204970 532170 205026 532226
rect 205094 532170 205150 532226
rect 205218 532170 205274 532226
rect 205342 532170 205398 532226
rect 204970 532046 205026 532102
rect 205094 532046 205150 532102
rect 205218 532046 205274 532102
rect 205342 532046 205398 532102
rect 204970 531922 205026 531978
rect 205094 531922 205150 531978
rect 205218 531922 205274 531978
rect 205342 531922 205398 531978
rect 204970 514294 205026 514350
rect 205094 514294 205150 514350
rect 205218 514294 205274 514350
rect 205342 514294 205398 514350
rect 204970 514170 205026 514226
rect 205094 514170 205150 514226
rect 205218 514170 205274 514226
rect 205342 514170 205398 514226
rect 204970 514046 205026 514102
rect 205094 514046 205150 514102
rect 205218 514046 205274 514102
rect 205342 514046 205398 514102
rect 204970 513922 205026 513978
rect 205094 513922 205150 513978
rect 205218 513922 205274 513978
rect 205342 513922 205398 513978
rect 204970 496294 205026 496350
rect 205094 496294 205150 496350
rect 205218 496294 205274 496350
rect 205342 496294 205398 496350
rect 204970 496170 205026 496226
rect 205094 496170 205150 496226
rect 205218 496170 205274 496226
rect 205342 496170 205398 496226
rect 204970 496046 205026 496102
rect 205094 496046 205150 496102
rect 205218 496046 205274 496102
rect 205342 496046 205398 496102
rect 204970 495922 205026 495978
rect 205094 495922 205150 495978
rect 205218 495922 205274 495978
rect 205342 495922 205398 495978
rect 204970 478294 205026 478350
rect 205094 478294 205150 478350
rect 205218 478294 205274 478350
rect 205342 478294 205398 478350
rect 204970 478170 205026 478226
rect 205094 478170 205150 478226
rect 205218 478170 205274 478226
rect 205342 478170 205398 478226
rect 204970 478046 205026 478102
rect 205094 478046 205150 478102
rect 205218 478046 205274 478102
rect 205342 478046 205398 478102
rect 204970 477922 205026 477978
rect 205094 477922 205150 477978
rect 205218 477922 205274 477978
rect 205342 477922 205398 477978
rect 204970 460294 205026 460350
rect 205094 460294 205150 460350
rect 205218 460294 205274 460350
rect 205342 460294 205398 460350
rect 204970 460170 205026 460226
rect 205094 460170 205150 460226
rect 205218 460170 205274 460226
rect 205342 460170 205398 460226
rect 204970 460046 205026 460102
rect 205094 460046 205150 460102
rect 205218 460046 205274 460102
rect 205342 460046 205398 460102
rect 204970 459922 205026 459978
rect 205094 459922 205150 459978
rect 205218 459922 205274 459978
rect 205342 459922 205398 459978
rect 204970 442294 205026 442350
rect 205094 442294 205150 442350
rect 205218 442294 205274 442350
rect 205342 442294 205398 442350
rect 204970 442170 205026 442226
rect 205094 442170 205150 442226
rect 205218 442170 205274 442226
rect 205342 442170 205398 442226
rect 204970 442046 205026 442102
rect 205094 442046 205150 442102
rect 205218 442046 205274 442102
rect 205342 442046 205398 442102
rect 204970 441922 205026 441978
rect 205094 441922 205150 441978
rect 205218 441922 205274 441978
rect 205342 441922 205398 441978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 219250 526294 219306 526350
rect 219374 526294 219430 526350
rect 219498 526294 219554 526350
rect 219622 526294 219678 526350
rect 219250 526170 219306 526226
rect 219374 526170 219430 526226
rect 219498 526170 219554 526226
rect 219622 526170 219678 526226
rect 219250 526046 219306 526102
rect 219374 526046 219430 526102
rect 219498 526046 219554 526102
rect 219622 526046 219678 526102
rect 219250 525922 219306 525978
rect 219374 525922 219430 525978
rect 219498 525922 219554 525978
rect 219622 525922 219678 525978
rect 219250 508294 219306 508350
rect 219374 508294 219430 508350
rect 219498 508294 219554 508350
rect 219622 508294 219678 508350
rect 219250 508170 219306 508226
rect 219374 508170 219430 508226
rect 219498 508170 219554 508226
rect 219622 508170 219678 508226
rect 219250 508046 219306 508102
rect 219374 508046 219430 508102
rect 219498 508046 219554 508102
rect 219622 508046 219678 508102
rect 219250 507922 219306 507978
rect 219374 507922 219430 507978
rect 219498 507922 219554 507978
rect 219622 507922 219678 507978
rect 219250 490294 219306 490350
rect 219374 490294 219430 490350
rect 219498 490294 219554 490350
rect 219622 490294 219678 490350
rect 219250 490170 219306 490226
rect 219374 490170 219430 490226
rect 219498 490170 219554 490226
rect 219622 490170 219678 490226
rect 219250 490046 219306 490102
rect 219374 490046 219430 490102
rect 219498 490046 219554 490102
rect 219622 490046 219678 490102
rect 219250 489922 219306 489978
rect 219374 489922 219430 489978
rect 219498 489922 219554 489978
rect 219622 489922 219678 489978
rect 219250 472294 219306 472350
rect 219374 472294 219430 472350
rect 219498 472294 219554 472350
rect 219622 472294 219678 472350
rect 219250 472170 219306 472226
rect 219374 472170 219430 472226
rect 219498 472170 219554 472226
rect 219622 472170 219678 472226
rect 219250 472046 219306 472102
rect 219374 472046 219430 472102
rect 219498 472046 219554 472102
rect 219622 472046 219678 472102
rect 219250 471922 219306 471978
rect 219374 471922 219430 471978
rect 219498 471922 219554 471978
rect 219622 471922 219678 471978
rect 219250 454294 219306 454350
rect 219374 454294 219430 454350
rect 219498 454294 219554 454350
rect 219622 454294 219678 454350
rect 219250 454170 219306 454226
rect 219374 454170 219430 454226
rect 219498 454170 219554 454226
rect 219622 454170 219678 454226
rect 219250 454046 219306 454102
rect 219374 454046 219430 454102
rect 219498 454046 219554 454102
rect 219622 454046 219678 454102
rect 219250 453922 219306 453978
rect 219374 453922 219430 453978
rect 219498 453922 219554 453978
rect 219622 453922 219678 453978
rect 218118 436261 218174 436317
rect 218242 436261 218298 436317
rect 218118 436137 218174 436193
rect 218242 436137 218298 436193
rect 218118 436013 218174 436069
rect 218242 436013 218298 436069
rect 187398 435889 187454 435945
rect 187522 435889 187578 435945
rect 219250 436322 219306 436378
rect 219374 436322 219430 436378
rect 219498 436322 219554 436378
rect 219622 436322 219678 436378
rect 219250 436198 219306 436254
rect 219374 436198 219430 436254
rect 219498 436198 219554 436254
rect 219622 436198 219678 436254
rect 219250 436074 219306 436130
rect 219374 436074 219430 436130
rect 219498 436074 219554 436130
rect 219622 436074 219678 436130
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 222970 514294 223026 514350
rect 223094 514294 223150 514350
rect 223218 514294 223274 514350
rect 223342 514294 223398 514350
rect 222970 514170 223026 514226
rect 223094 514170 223150 514226
rect 223218 514170 223274 514226
rect 223342 514170 223398 514226
rect 222970 514046 223026 514102
rect 223094 514046 223150 514102
rect 223218 514046 223274 514102
rect 223342 514046 223398 514102
rect 222970 513922 223026 513978
rect 223094 513922 223150 513978
rect 223218 513922 223274 513978
rect 223342 513922 223398 513978
rect 222970 496294 223026 496350
rect 223094 496294 223150 496350
rect 223218 496294 223274 496350
rect 223342 496294 223398 496350
rect 222970 496170 223026 496226
rect 223094 496170 223150 496226
rect 223218 496170 223274 496226
rect 223342 496170 223398 496226
rect 222970 496046 223026 496102
rect 223094 496046 223150 496102
rect 223218 496046 223274 496102
rect 223342 496046 223398 496102
rect 222970 495922 223026 495978
rect 223094 495922 223150 495978
rect 223218 495922 223274 495978
rect 223342 495922 223398 495978
rect 222970 478294 223026 478350
rect 223094 478294 223150 478350
rect 223218 478294 223274 478350
rect 223342 478294 223398 478350
rect 222970 478170 223026 478226
rect 223094 478170 223150 478226
rect 223218 478170 223274 478226
rect 223342 478170 223398 478226
rect 222970 478046 223026 478102
rect 223094 478046 223150 478102
rect 223218 478046 223274 478102
rect 223342 478046 223398 478102
rect 222970 477922 223026 477978
rect 223094 477922 223150 477978
rect 223218 477922 223274 477978
rect 223342 477922 223398 477978
rect 222970 460294 223026 460350
rect 223094 460294 223150 460350
rect 223218 460294 223274 460350
rect 223342 460294 223398 460350
rect 222970 460170 223026 460226
rect 223094 460170 223150 460226
rect 223218 460170 223274 460226
rect 223342 460170 223398 460226
rect 222970 460046 223026 460102
rect 223094 460046 223150 460102
rect 223218 460046 223274 460102
rect 223342 460046 223398 460102
rect 222970 459922 223026 459978
rect 223094 459922 223150 459978
rect 223218 459922 223274 459978
rect 223342 459922 223398 459978
rect 222970 442294 223026 442350
rect 223094 442294 223150 442350
rect 223218 442294 223274 442350
rect 223342 442294 223398 442350
rect 222970 442170 223026 442226
rect 223094 442170 223150 442226
rect 223218 442170 223274 442226
rect 223342 442170 223398 442226
rect 222970 442046 223026 442102
rect 223094 442046 223150 442102
rect 223218 442046 223274 442102
rect 223342 442046 223398 442102
rect 222970 441922 223026 441978
rect 223094 441922 223150 441978
rect 223218 441922 223274 441978
rect 223342 441922 223398 441978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 237250 526294 237306 526350
rect 237374 526294 237430 526350
rect 237498 526294 237554 526350
rect 237622 526294 237678 526350
rect 237250 526170 237306 526226
rect 237374 526170 237430 526226
rect 237498 526170 237554 526226
rect 237622 526170 237678 526226
rect 237250 526046 237306 526102
rect 237374 526046 237430 526102
rect 237498 526046 237554 526102
rect 237622 526046 237678 526102
rect 237250 525922 237306 525978
rect 237374 525922 237430 525978
rect 237498 525922 237554 525978
rect 237622 525922 237678 525978
rect 237250 508294 237306 508350
rect 237374 508294 237430 508350
rect 237498 508294 237554 508350
rect 237622 508294 237678 508350
rect 237250 508170 237306 508226
rect 237374 508170 237430 508226
rect 237498 508170 237554 508226
rect 237622 508170 237678 508226
rect 237250 508046 237306 508102
rect 237374 508046 237430 508102
rect 237498 508046 237554 508102
rect 237622 508046 237678 508102
rect 237250 507922 237306 507978
rect 237374 507922 237430 507978
rect 237498 507922 237554 507978
rect 237622 507922 237678 507978
rect 237250 490294 237306 490350
rect 237374 490294 237430 490350
rect 237498 490294 237554 490350
rect 237622 490294 237678 490350
rect 237250 490170 237306 490226
rect 237374 490170 237430 490226
rect 237498 490170 237554 490226
rect 237622 490170 237678 490226
rect 237250 490046 237306 490102
rect 237374 490046 237430 490102
rect 237498 490046 237554 490102
rect 237622 490046 237678 490102
rect 237250 489922 237306 489978
rect 237374 489922 237430 489978
rect 237498 489922 237554 489978
rect 237622 489922 237678 489978
rect 237250 472294 237306 472350
rect 237374 472294 237430 472350
rect 237498 472294 237554 472350
rect 237622 472294 237678 472350
rect 237250 472170 237306 472226
rect 237374 472170 237430 472226
rect 237498 472170 237554 472226
rect 237622 472170 237678 472226
rect 237250 472046 237306 472102
rect 237374 472046 237430 472102
rect 237498 472046 237554 472102
rect 237622 472046 237678 472102
rect 237250 471922 237306 471978
rect 237374 471922 237430 471978
rect 237498 471922 237554 471978
rect 237622 471922 237678 471978
rect 237250 454294 237306 454350
rect 237374 454294 237430 454350
rect 237498 454294 237554 454350
rect 237622 454294 237678 454350
rect 237250 454170 237306 454226
rect 237374 454170 237430 454226
rect 237498 454170 237554 454226
rect 237622 454170 237678 454226
rect 237250 454046 237306 454102
rect 237374 454046 237430 454102
rect 237498 454046 237554 454102
rect 237622 454046 237678 454102
rect 237250 453922 237306 453978
rect 237374 453922 237430 453978
rect 237498 453922 237554 453978
rect 237622 453922 237678 453978
rect 237250 436322 237306 436378
rect 237374 436322 237430 436378
rect 237498 436322 237554 436378
rect 237622 436322 237678 436378
rect 237250 436198 237306 436254
rect 237374 436198 237430 436254
rect 237498 436198 237554 436254
rect 237622 436198 237678 436254
rect 237250 436074 237306 436130
rect 237374 436074 237430 436130
rect 237498 436074 237554 436130
rect 237622 436074 237678 436130
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 240970 514294 241026 514350
rect 241094 514294 241150 514350
rect 241218 514294 241274 514350
rect 241342 514294 241398 514350
rect 240970 514170 241026 514226
rect 241094 514170 241150 514226
rect 241218 514170 241274 514226
rect 241342 514170 241398 514226
rect 240970 514046 241026 514102
rect 241094 514046 241150 514102
rect 241218 514046 241274 514102
rect 241342 514046 241398 514102
rect 240970 513922 241026 513978
rect 241094 513922 241150 513978
rect 241218 513922 241274 513978
rect 241342 513922 241398 513978
rect 240970 496294 241026 496350
rect 241094 496294 241150 496350
rect 241218 496294 241274 496350
rect 241342 496294 241398 496350
rect 240970 496170 241026 496226
rect 241094 496170 241150 496226
rect 241218 496170 241274 496226
rect 241342 496170 241398 496226
rect 240970 496046 241026 496102
rect 241094 496046 241150 496102
rect 241218 496046 241274 496102
rect 241342 496046 241398 496102
rect 240970 495922 241026 495978
rect 241094 495922 241150 495978
rect 241218 495922 241274 495978
rect 241342 495922 241398 495978
rect 240970 478294 241026 478350
rect 241094 478294 241150 478350
rect 241218 478294 241274 478350
rect 241342 478294 241398 478350
rect 240970 478170 241026 478226
rect 241094 478170 241150 478226
rect 241218 478170 241274 478226
rect 241342 478170 241398 478226
rect 240970 478046 241026 478102
rect 241094 478046 241150 478102
rect 241218 478046 241274 478102
rect 241342 478046 241398 478102
rect 240970 477922 241026 477978
rect 241094 477922 241150 477978
rect 241218 477922 241274 477978
rect 241342 477922 241398 477978
rect 240970 460294 241026 460350
rect 241094 460294 241150 460350
rect 241218 460294 241274 460350
rect 241342 460294 241398 460350
rect 240970 460170 241026 460226
rect 241094 460170 241150 460226
rect 241218 460170 241274 460226
rect 241342 460170 241398 460226
rect 240970 460046 241026 460102
rect 241094 460046 241150 460102
rect 241218 460046 241274 460102
rect 241342 460046 241398 460102
rect 240970 459922 241026 459978
rect 241094 459922 241150 459978
rect 241218 459922 241274 459978
rect 241342 459922 241398 459978
rect 240970 442294 241026 442350
rect 241094 442294 241150 442350
rect 241218 442294 241274 442350
rect 241342 442294 241398 442350
rect 240970 442170 241026 442226
rect 241094 442170 241150 442226
rect 241218 442170 241274 442226
rect 241342 442170 241398 442226
rect 240970 442046 241026 442102
rect 241094 442046 241150 442102
rect 241218 442046 241274 442102
rect 241342 442046 241398 442102
rect 240970 441922 241026 441978
rect 241094 441922 241150 441978
rect 241218 441922 241274 441978
rect 241342 441922 241398 441978
rect 255250 597156 255306 597212
rect 255374 597156 255430 597212
rect 255498 597156 255554 597212
rect 255622 597156 255678 597212
rect 255250 597032 255306 597088
rect 255374 597032 255430 597088
rect 255498 597032 255554 597088
rect 255622 597032 255678 597088
rect 255250 596908 255306 596964
rect 255374 596908 255430 596964
rect 255498 596908 255554 596964
rect 255622 596908 255678 596964
rect 255250 596784 255306 596840
rect 255374 596784 255430 596840
rect 255498 596784 255554 596840
rect 255622 596784 255678 596840
rect 255250 580294 255306 580350
rect 255374 580294 255430 580350
rect 255498 580294 255554 580350
rect 255622 580294 255678 580350
rect 255250 580170 255306 580226
rect 255374 580170 255430 580226
rect 255498 580170 255554 580226
rect 255622 580170 255678 580226
rect 255250 580046 255306 580102
rect 255374 580046 255430 580102
rect 255498 580046 255554 580102
rect 255622 580046 255678 580102
rect 255250 579922 255306 579978
rect 255374 579922 255430 579978
rect 255498 579922 255554 579978
rect 255622 579922 255678 579978
rect 255250 562294 255306 562350
rect 255374 562294 255430 562350
rect 255498 562294 255554 562350
rect 255622 562294 255678 562350
rect 255250 562170 255306 562226
rect 255374 562170 255430 562226
rect 255498 562170 255554 562226
rect 255622 562170 255678 562226
rect 255250 562046 255306 562102
rect 255374 562046 255430 562102
rect 255498 562046 255554 562102
rect 255622 562046 255678 562102
rect 255250 561922 255306 561978
rect 255374 561922 255430 561978
rect 255498 561922 255554 561978
rect 255622 561922 255678 561978
rect 255250 544294 255306 544350
rect 255374 544294 255430 544350
rect 255498 544294 255554 544350
rect 255622 544294 255678 544350
rect 255250 544170 255306 544226
rect 255374 544170 255430 544226
rect 255498 544170 255554 544226
rect 255622 544170 255678 544226
rect 255250 544046 255306 544102
rect 255374 544046 255430 544102
rect 255498 544046 255554 544102
rect 255622 544046 255678 544102
rect 255250 543922 255306 543978
rect 255374 543922 255430 543978
rect 255498 543922 255554 543978
rect 255622 543922 255678 543978
rect 255250 526294 255306 526350
rect 255374 526294 255430 526350
rect 255498 526294 255554 526350
rect 255622 526294 255678 526350
rect 255250 526170 255306 526226
rect 255374 526170 255430 526226
rect 255498 526170 255554 526226
rect 255622 526170 255678 526226
rect 255250 526046 255306 526102
rect 255374 526046 255430 526102
rect 255498 526046 255554 526102
rect 255622 526046 255678 526102
rect 255250 525922 255306 525978
rect 255374 525922 255430 525978
rect 255498 525922 255554 525978
rect 255622 525922 255678 525978
rect 255250 508294 255306 508350
rect 255374 508294 255430 508350
rect 255498 508294 255554 508350
rect 255622 508294 255678 508350
rect 255250 508170 255306 508226
rect 255374 508170 255430 508226
rect 255498 508170 255554 508226
rect 255622 508170 255678 508226
rect 255250 508046 255306 508102
rect 255374 508046 255430 508102
rect 255498 508046 255554 508102
rect 255622 508046 255678 508102
rect 255250 507922 255306 507978
rect 255374 507922 255430 507978
rect 255498 507922 255554 507978
rect 255622 507922 255678 507978
rect 255250 490294 255306 490350
rect 255374 490294 255430 490350
rect 255498 490294 255554 490350
rect 255622 490294 255678 490350
rect 255250 490170 255306 490226
rect 255374 490170 255430 490226
rect 255498 490170 255554 490226
rect 255622 490170 255678 490226
rect 255250 490046 255306 490102
rect 255374 490046 255430 490102
rect 255498 490046 255554 490102
rect 255622 490046 255678 490102
rect 255250 489922 255306 489978
rect 255374 489922 255430 489978
rect 255498 489922 255554 489978
rect 255622 489922 255678 489978
rect 255250 472294 255306 472350
rect 255374 472294 255430 472350
rect 255498 472294 255554 472350
rect 255622 472294 255678 472350
rect 255250 472170 255306 472226
rect 255374 472170 255430 472226
rect 255498 472170 255554 472226
rect 255622 472170 255678 472226
rect 255250 472046 255306 472102
rect 255374 472046 255430 472102
rect 255498 472046 255554 472102
rect 255622 472046 255678 472102
rect 255250 471922 255306 471978
rect 255374 471922 255430 471978
rect 255498 471922 255554 471978
rect 255622 471922 255678 471978
rect 255250 454294 255306 454350
rect 255374 454294 255430 454350
rect 255498 454294 255554 454350
rect 255622 454294 255678 454350
rect 255250 454170 255306 454226
rect 255374 454170 255430 454226
rect 255498 454170 255554 454226
rect 255622 454170 255678 454226
rect 255250 454046 255306 454102
rect 255374 454046 255430 454102
rect 255498 454046 255554 454102
rect 255622 454046 255678 454102
rect 255250 453922 255306 453978
rect 255374 453922 255430 453978
rect 255498 453922 255554 453978
rect 255622 453922 255678 453978
rect 248838 436261 248894 436317
rect 248962 436261 249018 436317
rect 248838 436137 248894 436193
rect 248962 436137 249018 436193
rect 248838 436013 248894 436069
rect 248962 436013 249018 436069
rect 218118 435889 218174 435945
rect 218242 435889 218298 435945
rect 255250 436322 255306 436378
rect 255374 436322 255430 436378
rect 255498 436322 255554 436378
rect 255622 436322 255678 436378
rect 255250 436198 255306 436254
rect 255374 436198 255430 436254
rect 255498 436198 255554 436254
rect 255622 436198 255678 436254
rect 255250 436074 255306 436130
rect 255374 436074 255430 436130
rect 255498 436074 255554 436130
rect 255622 436074 255678 436130
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 258970 514294 259026 514350
rect 259094 514294 259150 514350
rect 259218 514294 259274 514350
rect 259342 514294 259398 514350
rect 258970 514170 259026 514226
rect 259094 514170 259150 514226
rect 259218 514170 259274 514226
rect 259342 514170 259398 514226
rect 258970 514046 259026 514102
rect 259094 514046 259150 514102
rect 259218 514046 259274 514102
rect 259342 514046 259398 514102
rect 258970 513922 259026 513978
rect 259094 513922 259150 513978
rect 259218 513922 259274 513978
rect 259342 513922 259398 513978
rect 258970 496294 259026 496350
rect 259094 496294 259150 496350
rect 259218 496294 259274 496350
rect 259342 496294 259398 496350
rect 258970 496170 259026 496226
rect 259094 496170 259150 496226
rect 259218 496170 259274 496226
rect 259342 496170 259398 496226
rect 258970 496046 259026 496102
rect 259094 496046 259150 496102
rect 259218 496046 259274 496102
rect 259342 496046 259398 496102
rect 258970 495922 259026 495978
rect 259094 495922 259150 495978
rect 259218 495922 259274 495978
rect 259342 495922 259398 495978
rect 258970 478294 259026 478350
rect 259094 478294 259150 478350
rect 259218 478294 259274 478350
rect 259342 478294 259398 478350
rect 258970 478170 259026 478226
rect 259094 478170 259150 478226
rect 259218 478170 259274 478226
rect 259342 478170 259398 478226
rect 258970 478046 259026 478102
rect 259094 478046 259150 478102
rect 259218 478046 259274 478102
rect 259342 478046 259398 478102
rect 258970 477922 259026 477978
rect 259094 477922 259150 477978
rect 259218 477922 259274 477978
rect 259342 477922 259398 477978
rect 258970 460294 259026 460350
rect 259094 460294 259150 460350
rect 259218 460294 259274 460350
rect 259342 460294 259398 460350
rect 258970 460170 259026 460226
rect 259094 460170 259150 460226
rect 259218 460170 259274 460226
rect 259342 460170 259398 460226
rect 258970 460046 259026 460102
rect 259094 460046 259150 460102
rect 259218 460046 259274 460102
rect 259342 460046 259398 460102
rect 258970 459922 259026 459978
rect 259094 459922 259150 459978
rect 259218 459922 259274 459978
rect 259342 459922 259398 459978
rect 258970 442294 259026 442350
rect 259094 442294 259150 442350
rect 259218 442294 259274 442350
rect 259342 442294 259398 442350
rect 258970 442170 259026 442226
rect 259094 442170 259150 442226
rect 259218 442170 259274 442226
rect 259342 442170 259398 442226
rect 258970 442046 259026 442102
rect 259094 442046 259150 442102
rect 259218 442046 259274 442102
rect 259342 442046 259398 442102
rect 258970 441922 259026 441978
rect 259094 441922 259150 441978
rect 259218 441922 259274 441978
rect 259342 441922 259398 441978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 273250 526294 273306 526350
rect 273374 526294 273430 526350
rect 273498 526294 273554 526350
rect 273622 526294 273678 526350
rect 273250 526170 273306 526226
rect 273374 526170 273430 526226
rect 273498 526170 273554 526226
rect 273622 526170 273678 526226
rect 273250 526046 273306 526102
rect 273374 526046 273430 526102
rect 273498 526046 273554 526102
rect 273622 526046 273678 526102
rect 273250 525922 273306 525978
rect 273374 525922 273430 525978
rect 273498 525922 273554 525978
rect 273622 525922 273678 525978
rect 273250 508294 273306 508350
rect 273374 508294 273430 508350
rect 273498 508294 273554 508350
rect 273622 508294 273678 508350
rect 273250 508170 273306 508226
rect 273374 508170 273430 508226
rect 273498 508170 273554 508226
rect 273622 508170 273678 508226
rect 273250 508046 273306 508102
rect 273374 508046 273430 508102
rect 273498 508046 273554 508102
rect 273622 508046 273678 508102
rect 273250 507922 273306 507978
rect 273374 507922 273430 507978
rect 273498 507922 273554 507978
rect 273622 507922 273678 507978
rect 273250 490294 273306 490350
rect 273374 490294 273430 490350
rect 273498 490294 273554 490350
rect 273622 490294 273678 490350
rect 273250 490170 273306 490226
rect 273374 490170 273430 490226
rect 273498 490170 273554 490226
rect 273622 490170 273678 490226
rect 273250 490046 273306 490102
rect 273374 490046 273430 490102
rect 273498 490046 273554 490102
rect 273622 490046 273678 490102
rect 273250 489922 273306 489978
rect 273374 489922 273430 489978
rect 273498 489922 273554 489978
rect 273622 489922 273678 489978
rect 273250 472294 273306 472350
rect 273374 472294 273430 472350
rect 273498 472294 273554 472350
rect 273622 472294 273678 472350
rect 273250 472170 273306 472226
rect 273374 472170 273430 472226
rect 273498 472170 273554 472226
rect 273622 472170 273678 472226
rect 273250 472046 273306 472102
rect 273374 472046 273430 472102
rect 273498 472046 273554 472102
rect 273622 472046 273678 472102
rect 273250 471922 273306 471978
rect 273374 471922 273430 471978
rect 273498 471922 273554 471978
rect 273622 471922 273678 471978
rect 273250 454294 273306 454350
rect 273374 454294 273430 454350
rect 273498 454294 273554 454350
rect 273622 454294 273678 454350
rect 273250 454170 273306 454226
rect 273374 454170 273430 454226
rect 273498 454170 273554 454226
rect 273622 454170 273678 454226
rect 273250 454046 273306 454102
rect 273374 454046 273430 454102
rect 273498 454046 273554 454102
rect 273622 454046 273678 454102
rect 273250 453922 273306 453978
rect 273374 453922 273430 453978
rect 273498 453922 273554 453978
rect 273622 453922 273678 453978
rect 273250 436322 273306 436378
rect 273374 436322 273430 436378
rect 273498 436322 273554 436378
rect 273622 436322 273678 436378
rect 273250 436198 273306 436254
rect 273374 436198 273430 436254
rect 273498 436198 273554 436254
rect 273622 436198 273678 436254
rect 273250 436074 273306 436130
rect 273374 436074 273430 436130
rect 273498 436074 273554 436130
rect 273622 436074 273678 436130
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 276970 514294 277026 514350
rect 277094 514294 277150 514350
rect 277218 514294 277274 514350
rect 277342 514294 277398 514350
rect 276970 514170 277026 514226
rect 277094 514170 277150 514226
rect 277218 514170 277274 514226
rect 277342 514170 277398 514226
rect 276970 514046 277026 514102
rect 277094 514046 277150 514102
rect 277218 514046 277274 514102
rect 277342 514046 277398 514102
rect 276970 513922 277026 513978
rect 277094 513922 277150 513978
rect 277218 513922 277274 513978
rect 277342 513922 277398 513978
rect 276970 496294 277026 496350
rect 277094 496294 277150 496350
rect 277218 496294 277274 496350
rect 277342 496294 277398 496350
rect 276970 496170 277026 496226
rect 277094 496170 277150 496226
rect 277218 496170 277274 496226
rect 277342 496170 277398 496226
rect 276970 496046 277026 496102
rect 277094 496046 277150 496102
rect 277218 496046 277274 496102
rect 277342 496046 277398 496102
rect 276970 495922 277026 495978
rect 277094 495922 277150 495978
rect 277218 495922 277274 495978
rect 277342 495922 277398 495978
rect 276970 478294 277026 478350
rect 277094 478294 277150 478350
rect 277218 478294 277274 478350
rect 277342 478294 277398 478350
rect 276970 478170 277026 478226
rect 277094 478170 277150 478226
rect 277218 478170 277274 478226
rect 277342 478170 277398 478226
rect 276970 478046 277026 478102
rect 277094 478046 277150 478102
rect 277218 478046 277274 478102
rect 277342 478046 277398 478102
rect 276970 477922 277026 477978
rect 277094 477922 277150 477978
rect 277218 477922 277274 477978
rect 277342 477922 277398 477978
rect 276970 460294 277026 460350
rect 277094 460294 277150 460350
rect 277218 460294 277274 460350
rect 277342 460294 277398 460350
rect 276970 460170 277026 460226
rect 277094 460170 277150 460226
rect 277218 460170 277274 460226
rect 277342 460170 277398 460226
rect 276970 460046 277026 460102
rect 277094 460046 277150 460102
rect 277218 460046 277274 460102
rect 277342 460046 277398 460102
rect 276970 459922 277026 459978
rect 277094 459922 277150 459978
rect 277218 459922 277274 459978
rect 277342 459922 277398 459978
rect 276970 442294 277026 442350
rect 277094 442294 277150 442350
rect 277218 442294 277274 442350
rect 277342 442294 277398 442350
rect 276970 442170 277026 442226
rect 277094 442170 277150 442226
rect 277218 442170 277274 442226
rect 277342 442170 277398 442226
rect 276970 442046 277026 442102
rect 277094 442046 277150 442102
rect 277218 442046 277274 442102
rect 277342 442046 277398 442102
rect 276970 441922 277026 441978
rect 277094 441922 277150 441978
rect 277218 441922 277274 441978
rect 277342 441922 277398 441978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 291250 526294 291306 526350
rect 291374 526294 291430 526350
rect 291498 526294 291554 526350
rect 291622 526294 291678 526350
rect 291250 526170 291306 526226
rect 291374 526170 291430 526226
rect 291498 526170 291554 526226
rect 291622 526170 291678 526226
rect 291250 526046 291306 526102
rect 291374 526046 291430 526102
rect 291498 526046 291554 526102
rect 291622 526046 291678 526102
rect 291250 525922 291306 525978
rect 291374 525922 291430 525978
rect 291498 525922 291554 525978
rect 291622 525922 291678 525978
rect 291250 508294 291306 508350
rect 291374 508294 291430 508350
rect 291498 508294 291554 508350
rect 291622 508294 291678 508350
rect 291250 508170 291306 508226
rect 291374 508170 291430 508226
rect 291498 508170 291554 508226
rect 291622 508170 291678 508226
rect 291250 508046 291306 508102
rect 291374 508046 291430 508102
rect 291498 508046 291554 508102
rect 291622 508046 291678 508102
rect 291250 507922 291306 507978
rect 291374 507922 291430 507978
rect 291498 507922 291554 507978
rect 291622 507922 291678 507978
rect 291250 490294 291306 490350
rect 291374 490294 291430 490350
rect 291498 490294 291554 490350
rect 291622 490294 291678 490350
rect 291250 490170 291306 490226
rect 291374 490170 291430 490226
rect 291498 490170 291554 490226
rect 291622 490170 291678 490226
rect 291250 490046 291306 490102
rect 291374 490046 291430 490102
rect 291498 490046 291554 490102
rect 291622 490046 291678 490102
rect 291250 489922 291306 489978
rect 291374 489922 291430 489978
rect 291498 489922 291554 489978
rect 291622 489922 291678 489978
rect 291250 472294 291306 472350
rect 291374 472294 291430 472350
rect 291498 472294 291554 472350
rect 291622 472294 291678 472350
rect 291250 472170 291306 472226
rect 291374 472170 291430 472226
rect 291498 472170 291554 472226
rect 291622 472170 291678 472226
rect 291250 472046 291306 472102
rect 291374 472046 291430 472102
rect 291498 472046 291554 472102
rect 291622 472046 291678 472102
rect 291250 471922 291306 471978
rect 291374 471922 291430 471978
rect 291498 471922 291554 471978
rect 291622 471922 291678 471978
rect 291250 454294 291306 454350
rect 291374 454294 291430 454350
rect 291498 454294 291554 454350
rect 291622 454294 291678 454350
rect 291250 454170 291306 454226
rect 291374 454170 291430 454226
rect 291498 454170 291554 454226
rect 291622 454170 291678 454226
rect 291250 454046 291306 454102
rect 291374 454046 291430 454102
rect 291498 454046 291554 454102
rect 291622 454046 291678 454102
rect 291250 453922 291306 453978
rect 291374 453922 291430 453978
rect 291498 453922 291554 453978
rect 291622 453922 291678 453978
rect 279558 436261 279614 436317
rect 279682 436261 279738 436317
rect 279558 436137 279614 436193
rect 279682 436137 279738 436193
rect 279558 436013 279614 436069
rect 279682 436013 279738 436069
rect 248838 435889 248894 435945
rect 248962 435889 249018 435945
rect 294970 598116 295026 598172
rect 295094 598116 295150 598172
rect 295218 598116 295274 598172
rect 295342 598116 295398 598172
rect 294970 597992 295026 598048
rect 295094 597992 295150 598048
rect 295218 597992 295274 598048
rect 295342 597992 295398 598048
rect 294970 597868 295026 597924
rect 295094 597868 295150 597924
rect 295218 597868 295274 597924
rect 295342 597868 295398 597924
rect 294970 597744 295026 597800
rect 295094 597744 295150 597800
rect 295218 597744 295274 597800
rect 295342 597744 295398 597800
rect 294970 586294 295026 586350
rect 295094 586294 295150 586350
rect 295218 586294 295274 586350
rect 295342 586294 295398 586350
rect 294970 586170 295026 586226
rect 295094 586170 295150 586226
rect 295218 586170 295274 586226
rect 295342 586170 295398 586226
rect 294970 586046 295026 586102
rect 295094 586046 295150 586102
rect 295218 586046 295274 586102
rect 295342 586046 295398 586102
rect 294970 585922 295026 585978
rect 295094 585922 295150 585978
rect 295218 585922 295274 585978
rect 295342 585922 295398 585978
rect 294970 568294 295026 568350
rect 295094 568294 295150 568350
rect 295218 568294 295274 568350
rect 295342 568294 295398 568350
rect 294970 568170 295026 568226
rect 295094 568170 295150 568226
rect 295218 568170 295274 568226
rect 295342 568170 295398 568226
rect 294970 568046 295026 568102
rect 295094 568046 295150 568102
rect 295218 568046 295274 568102
rect 295342 568046 295398 568102
rect 294970 567922 295026 567978
rect 295094 567922 295150 567978
rect 295218 567922 295274 567978
rect 295342 567922 295398 567978
rect 294970 550294 295026 550350
rect 295094 550294 295150 550350
rect 295218 550294 295274 550350
rect 295342 550294 295398 550350
rect 294970 550170 295026 550226
rect 295094 550170 295150 550226
rect 295218 550170 295274 550226
rect 295342 550170 295398 550226
rect 294970 550046 295026 550102
rect 295094 550046 295150 550102
rect 295218 550046 295274 550102
rect 295342 550046 295398 550102
rect 294970 549922 295026 549978
rect 295094 549922 295150 549978
rect 295218 549922 295274 549978
rect 295342 549922 295398 549978
rect 294970 532294 295026 532350
rect 295094 532294 295150 532350
rect 295218 532294 295274 532350
rect 295342 532294 295398 532350
rect 294970 532170 295026 532226
rect 295094 532170 295150 532226
rect 295218 532170 295274 532226
rect 295342 532170 295398 532226
rect 294970 532046 295026 532102
rect 295094 532046 295150 532102
rect 295218 532046 295274 532102
rect 295342 532046 295398 532102
rect 294970 531922 295026 531978
rect 295094 531922 295150 531978
rect 295218 531922 295274 531978
rect 295342 531922 295398 531978
rect 294970 514294 295026 514350
rect 295094 514294 295150 514350
rect 295218 514294 295274 514350
rect 295342 514294 295398 514350
rect 294970 514170 295026 514226
rect 295094 514170 295150 514226
rect 295218 514170 295274 514226
rect 295342 514170 295398 514226
rect 294970 514046 295026 514102
rect 295094 514046 295150 514102
rect 295218 514046 295274 514102
rect 295342 514046 295398 514102
rect 294970 513922 295026 513978
rect 295094 513922 295150 513978
rect 295218 513922 295274 513978
rect 295342 513922 295398 513978
rect 294970 496294 295026 496350
rect 295094 496294 295150 496350
rect 295218 496294 295274 496350
rect 295342 496294 295398 496350
rect 294970 496170 295026 496226
rect 295094 496170 295150 496226
rect 295218 496170 295274 496226
rect 295342 496170 295398 496226
rect 294970 496046 295026 496102
rect 295094 496046 295150 496102
rect 295218 496046 295274 496102
rect 295342 496046 295398 496102
rect 294970 495922 295026 495978
rect 295094 495922 295150 495978
rect 295218 495922 295274 495978
rect 295342 495922 295398 495978
rect 294970 478294 295026 478350
rect 295094 478294 295150 478350
rect 295218 478294 295274 478350
rect 295342 478294 295398 478350
rect 294970 478170 295026 478226
rect 295094 478170 295150 478226
rect 295218 478170 295274 478226
rect 295342 478170 295398 478226
rect 294970 478046 295026 478102
rect 295094 478046 295150 478102
rect 295218 478046 295274 478102
rect 295342 478046 295398 478102
rect 294970 477922 295026 477978
rect 295094 477922 295150 477978
rect 295218 477922 295274 477978
rect 295342 477922 295398 477978
rect 294970 460294 295026 460350
rect 295094 460294 295150 460350
rect 295218 460294 295274 460350
rect 295342 460294 295398 460350
rect 294970 460170 295026 460226
rect 295094 460170 295150 460226
rect 295218 460170 295274 460226
rect 295342 460170 295398 460226
rect 294970 460046 295026 460102
rect 295094 460046 295150 460102
rect 295218 460046 295274 460102
rect 295342 460046 295398 460102
rect 294970 459922 295026 459978
rect 295094 459922 295150 459978
rect 295218 459922 295274 459978
rect 295342 459922 295398 459978
rect 294970 442294 295026 442350
rect 295094 442294 295150 442350
rect 295218 442294 295274 442350
rect 295342 442294 295398 442350
rect 294970 442170 295026 442226
rect 295094 442170 295150 442226
rect 295218 442170 295274 442226
rect 295342 442170 295398 442226
rect 294970 442046 295026 442102
rect 295094 442046 295150 442102
rect 295218 442046 295274 442102
rect 295342 442046 295398 442102
rect 294970 441922 295026 441978
rect 295094 441922 295150 441978
rect 295218 441922 295274 441978
rect 295342 441922 295398 441978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 309250 526294 309306 526350
rect 309374 526294 309430 526350
rect 309498 526294 309554 526350
rect 309622 526294 309678 526350
rect 309250 526170 309306 526226
rect 309374 526170 309430 526226
rect 309498 526170 309554 526226
rect 309622 526170 309678 526226
rect 309250 526046 309306 526102
rect 309374 526046 309430 526102
rect 309498 526046 309554 526102
rect 309622 526046 309678 526102
rect 309250 525922 309306 525978
rect 309374 525922 309430 525978
rect 309498 525922 309554 525978
rect 309622 525922 309678 525978
rect 309250 508294 309306 508350
rect 309374 508294 309430 508350
rect 309498 508294 309554 508350
rect 309622 508294 309678 508350
rect 309250 508170 309306 508226
rect 309374 508170 309430 508226
rect 309498 508170 309554 508226
rect 309622 508170 309678 508226
rect 309250 508046 309306 508102
rect 309374 508046 309430 508102
rect 309498 508046 309554 508102
rect 309622 508046 309678 508102
rect 309250 507922 309306 507978
rect 309374 507922 309430 507978
rect 309498 507922 309554 507978
rect 309622 507922 309678 507978
rect 309250 490294 309306 490350
rect 309374 490294 309430 490350
rect 309498 490294 309554 490350
rect 309622 490294 309678 490350
rect 309250 490170 309306 490226
rect 309374 490170 309430 490226
rect 309498 490170 309554 490226
rect 309622 490170 309678 490226
rect 309250 490046 309306 490102
rect 309374 490046 309430 490102
rect 309498 490046 309554 490102
rect 309622 490046 309678 490102
rect 309250 489922 309306 489978
rect 309374 489922 309430 489978
rect 309498 489922 309554 489978
rect 309622 489922 309678 489978
rect 309250 472294 309306 472350
rect 309374 472294 309430 472350
rect 309498 472294 309554 472350
rect 309622 472294 309678 472350
rect 309250 472170 309306 472226
rect 309374 472170 309430 472226
rect 309498 472170 309554 472226
rect 309622 472170 309678 472226
rect 309250 472046 309306 472102
rect 309374 472046 309430 472102
rect 309498 472046 309554 472102
rect 309622 472046 309678 472102
rect 309250 471922 309306 471978
rect 309374 471922 309430 471978
rect 309498 471922 309554 471978
rect 309622 471922 309678 471978
rect 309250 454294 309306 454350
rect 309374 454294 309430 454350
rect 309498 454294 309554 454350
rect 309622 454294 309678 454350
rect 309250 454170 309306 454226
rect 309374 454170 309430 454226
rect 309498 454170 309554 454226
rect 309622 454170 309678 454226
rect 309250 454046 309306 454102
rect 309374 454046 309430 454102
rect 309498 454046 309554 454102
rect 309622 454046 309678 454102
rect 309250 453922 309306 453978
rect 309374 453922 309430 453978
rect 309498 453922 309554 453978
rect 309622 453922 309678 453978
rect 291250 436322 291306 436378
rect 291374 436322 291430 436378
rect 291498 436322 291554 436378
rect 291622 436322 291678 436378
rect 291250 436198 291306 436254
rect 291374 436198 291430 436254
rect 291498 436198 291554 436254
rect 291622 436198 291678 436254
rect 291250 436074 291306 436130
rect 291374 436074 291430 436130
rect 291498 436074 291554 436130
rect 291622 436074 291678 436130
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 312970 514294 313026 514350
rect 313094 514294 313150 514350
rect 313218 514294 313274 514350
rect 313342 514294 313398 514350
rect 312970 514170 313026 514226
rect 313094 514170 313150 514226
rect 313218 514170 313274 514226
rect 313342 514170 313398 514226
rect 312970 514046 313026 514102
rect 313094 514046 313150 514102
rect 313218 514046 313274 514102
rect 313342 514046 313398 514102
rect 312970 513922 313026 513978
rect 313094 513922 313150 513978
rect 313218 513922 313274 513978
rect 313342 513922 313398 513978
rect 312970 496294 313026 496350
rect 313094 496294 313150 496350
rect 313218 496294 313274 496350
rect 313342 496294 313398 496350
rect 312970 496170 313026 496226
rect 313094 496170 313150 496226
rect 313218 496170 313274 496226
rect 313342 496170 313398 496226
rect 312970 496046 313026 496102
rect 313094 496046 313150 496102
rect 313218 496046 313274 496102
rect 313342 496046 313398 496102
rect 312970 495922 313026 495978
rect 313094 495922 313150 495978
rect 313218 495922 313274 495978
rect 313342 495922 313398 495978
rect 312970 478294 313026 478350
rect 313094 478294 313150 478350
rect 313218 478294 313274 478350
rect 313342 478294 313398 478350
rect 312970 478170 313026 478226
rect 313094 478170 313150 478226
rect 313218 478170 313274 478226
rect 313342 478170 313398 478226
rect 312970 478046 313026 478102
rect 313094 478046 313150 478102
rect 313218 478046 313274 478102
rect 313342 478046 313398 478102
rect 312970 477922 313026 477978
rect 313094 477922 313150 477978
rect 313218 477922 313274 477978
rect 313342 477922 313398 477978
rect 312970 460294 313026 460350
rect 313094 460294 313150 460350
rect 313218 460294 313274 460350
rect 313342 460294 313398 460350
rect 312970 460170 313026 460226
rect 313094 460170 313150 460226
rect 313218 460170 313274 460226
rect 313342 460170 313398 460226
rect 312970 460046 313026 460102
rect 313094 460046 313150 460102
rect 313218 460046 313274 460102
rect 313342 460046 313398 460102
rect 312970 459922 313026 459978
rect 313094 459922 313150 459978
rect 313218 459922 313274 459978
rect 313342 459922 313398 459978
rect 312970 442294 313026 442350
rect 313094 442294 313150 442350
rect 313218 442294 313274 442350
rect 313342 442294 313398 442350
rect 312970 442170 313026 442226
rect 313094 442170 313150 442226
rect 313218 442170 313274 442226
rect 313342 442170 313398 442226
rect 312970 442046 313026 442102
rect 313094 442046 313150 442102
rect 313218 442046 313274 442102
rect 313342 442046 313398 442102
rect 312970 441922 313026 441978
rect 313094 441922 313150 441978
rect 313218 441922 313274 441978
rect 313342 441922 313398 441978
rect 309250 436322 309306 436378
rect 309374 436322 309430 436378
rect 309498 436322 309554 436378
rect 309622 436322 309678 436378
rect 309250 436198 309306 436254
rect 309374 436198 309430 436254
rect 309498 436198 309554 436254
rect 309622 436198 309678 436254
rect 309250 436074 309306 436130
rect 309374 436074 309430 436130
rect 309498 436074 309554 436130
rect 309622 436074 309678 436130
rect 310278 436261 310334 436317
rect 310402 436261 310458 436317
rect 310278 436137 310334 436193
rect 310402 436137 310458 436193
rect 310278 436013 310334 436069
rect 310402 436013 310458 436069
rect 279558 435889 279614 435945
rect 279682 435889 279738 435945
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 327250 526294 327306 526350
rect 327374 526294 327430 526350
rect 327498 526294 327554 526350
rect 327622 526294 327678 526350
rect 327250 526170 327306 526226
rect 327374 526170 327430 526226
rect 327498 526170 327554 526226
rect 327622 526170 327678 526226
rect 327250 526046 327306 526102
rect 327374 526046 327430 526102
rect 327498 526046 327554 526102
rect 327622 526046 327678 526102
rect 327250 525922 327306 525978
rect 327374 525922 327430 525978
rect 327498 525922 327554 525978
rect 327622 525922 327678 525978
rect 327250 508294 327306 508350
rect 327374 508294 327430 508350
rect 327498 508294 327554 508350
rect 327622 508294 327678 508350
rect 327250 508170 327306 508226
rect 327374 508170 327430 508226
rect 327498 508170 327554 508226
rect 327622 508170 327678 508226
rect 327250 508046 327306 508102
rect 327374 508046 327430 508102
rect 327498 508046 327554 508102
rect 327622 508046 327678 508102
rect 327250 507922 327306 507978
rect 327374 507922 327430 507978
rect 327498 507922 327554 507978
rect 327622 507922 327678 507978
rect 327250 490294 327306 490350
rect 327374 490294 327430 490350
rect 327498 490294 327554 490350
rect 327622 490294 327678 490350
rect 327250 490170 327306 490226
rect 327374 490170 327430 490226
rect 327498 490170 327554 490226
rect 327622 490170 327678 490226
rect 327250 490046 327306 490102
rect 327374 490046 327430 490102
rect 327498 490046 327554 490102
rect 327622 490046 327678 490102
rect 327250 489922 327306 489978
rect 327374 489922 327430 489978
rect 327498 489922 327554 489978
rect 327622 489922 327678 489978
rect 327250 472294 327306 472350
rect 327374 472294 327430 472350
rect 327498 472294 327554 472350
rect 327622 472294 327678 472350
rect 327250 472170 327306 472226
rect 327374 472170 327430 472226
rect 327498 472170 327554 472226
rect 327622 472170 327678 472226
rect 327250 472046 327306 472102
rect 327374 472046 327430 472102
rect 327498 472046 327554 472102
rect 327622 472046 327678 472102
rect 327250 471922 327306 471978
rect 327374 471922 327430 471978
rect 327498 471922 327554 471978
rect 327622 471922 327678 471978
rect 327250 454294 327306 454350
rect 327374 454294 327430 454350
rect 327498 454294 327554 454350
rect 327622 454294 327678 454350
rect 327250 454170 327306 454226
rect 327374 454170 327430 454226
rect 327498 454170 327554 454226
rect 327622 454170 327678 454226
rect 327250 454046 327306 454102
rect 327374 454046 327430 454102
rect 327498 454046 327554 454102
rect 327622 454046 327678 454102
rect 327250 453922 327306 453978
rect 327374 453922 327430 453978
rect 327498 453922 327554 453978
rect 327622 453922 327678 453978
rect 327250 436322 327306 436378
rect 327374 436322 327430 436378
rect 327498 436322 327554 436378
rect 327622 436322 327678 436378
rect 327250 436198 327306 436254
rect 327374 436198 327430 436254
rect 327498 436198 327554 436254
rect 327622 436198 327678 436254
rect 327250 436074 327306 436130
rect 327374 436074 327430 436130
rect 327498 436074 327554 436130
rect 327622 436074 327678 436130
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 330970 514294 331026 514350
rect 331094 514294 331150 514350
rect 331218 514294 331274 514350
rect 331342 514294 331398 514350
rect 330970 514170 331026 514226
rect 331094 514170 331150 514226
rect 331218 514170 331274 514226
rect 331342 514170 331398 514226
rect 330970 514046 331026 514102
rect 331094 514046 331150 514102
rect 331218 514046 331274 514102
rect 331342 514046 331398 514102
rect 330970 513922 331026 513978
rect 331094 513922 331150 513978
rect 331218 513922 331274 513978
rect 331342 513922 331398 513978
rect 330970 496294 331026 496350
rect 331094 496294 331150 496350
rect 331218 496294 331274 496350
rect 331342 496294 331398 496350
rect 330970 496170 331026 496226
rect 331094 496170 331150 496226
rect 331218 496170 331274 496226
rect 331342 496170 331398 496226
rect 330970 496046 331026 496102
rect 331094 496046 331150 496102
rect 331218 496046 331274 496102
rect 331342 496046 331398 496102
rect 330970 495922 331026 495978
rect 331094 495922 331150 495978
rect 331218 495922 331274 495978
rect 331342 495922 331398 495978
rect 330970 478294 331026 478350
rect 331094 478294 331150 478350
rect 331218 478294 331274 478350
rect 331342 478294 331398 478350
rect 330970 478170 331026 478226
rect 331094 478170 331150 478226
rect 331218 478170 331274 478226
rect 331342 478170 331398 478226
rect 330970 478046 331026 478102
rect 331094 478046 331150 478102
rect 331218 478046 331274 478102
rect 331342 478046 331398 478102
rect 330970 477922 331026 477978
rect 331094 477922 331150 477978
rect 331218 477922 331274 477978
rect 331342 477922 331398 477978
rect 330970 460294 331026 460350
rect 331094 460294 331150 460350
rect 331218 460294 331274 460350
rect 331342 460294 331398 460350
rect 330970 460170 331026 460226
rect 331094 460170 331150 460226
rect 331218 460170 331274 460226
rect 331342 460170 331398 460226
rect 330970 460046 331026 460102
rect 331094 460046 331150 460102
rect 331218 460046 331274 460102
rect 331342 460046 331398 460102
rect 330970 459922 331026 459978
rect 331094 459922 331150 459978
rect 331218 459922 331274 459978
rect 331342 459922 331398 459978
rect 330970 442294 331026 442350
rect 331094 442294 331150 442350
rect 331218 442294 331274 442350
rect 331342 442294 331398 442350
rect 330970 442170 331026 442226
rect 331094 442170 331150 442226
rect 331218 442170 331274 442226
rect 331342 442170 331398 442226
rect 330970 442046 331026 442102
rect 331094 442046 331150 442102
rect 331218 442046 331274 442102
rect 331342 442046 331398 442102
rect 330970 441922 331026 441978
rect 331094 441922 331150 441978
rect 331218 441922 331274 441978
rect 331342 441922 331398 441978
rect 345250 597156 345306 597212
rect 345374 597156 345430 597212
rect 345498 597156 345554 597212
rect 345622 597156 345678 597212
rect 345250 597032 345306 597088
rect 345374 597032 345430 597088
rect 345498 597032 345554 597088
rect 345622 597032 345678 597088
rect 345250 596908 345306 596964
rect 345374 596908 345430 596964
rect 345498 596908 345554 596964
rect 345622 596908 345678 596964
rect 345250 596784 345306 596840
rect 345374 596784 345430 596840
rect 345498 596784 345554 596840
rect 345622 596784 345678 596840
rect 345250 580294 345306 580350
rect 345374 580294 345430 580350
rect 345498 580294 345554 580350
rect 345622 580294 345678 580350
rect 345250 580170 345306 580226
rect 345374 580170 345430 580226
rect 345498 580170 345554 580226
rect 345622 580170 345678 580226
rect 345250 580046 345306 580102
rect 345374 580046 345430 580102
rect 345498 580046 345554 580102
rect 345622 580046 345678 580102
rect 345250 579922 345306 579978
rect 345374 579922 345430 579978
rect 345498 579922 345554 579978
rect 345622 579922 345678 579978
rect 345250 562294 345306 562350
rect 345374 562294 345430 562350
rect 345498 562294 345554 562350
rect 345622 562294 345678 562350
rect 345250 562170 345306 562226
rect 345374 562170 345430 562226
rect 345498 562170 345554 562226
rect 345622 562170 345678 562226
rect 345250 562046 345306 562102
rect 345374 562046 345430 562102
rect 345498 562046 345554 562102
rect 345622 562046 345678 562102
rect 345250 561922 345306 561978
rect 345374 561922 345430 561978
rect 345498 561922 345554 561978
rect 345622 561922 345678 561978
rect 345250 544294 345306 544350
rect 345374 544294 345430 544350
rect 345498 544294 345554 544350
rect 345622 544294 345678 544350
rect 345250 544170 345306 544226
rect 345374 544170 345430 544226
rect 345498 544170 345554 544226
rect 345622 544170 345678 544226
rect 345250 544046 345306 544102
rect 345374 544046 345430 544102
rect 345498 544046 345554 544102
rect 345622 544046 345678 544102
rect 345250 543922 345306 543978
rect 345374 543922 345430 543978
rect 345498 543922 345554 543978
rect 345622 543922 345678 543978
rect 345250 526294 345306 526350
rect 345374 526294 345430 526350
rect 345498 526294 345554 526350
rect 345622 526294 345678 526350
rect 345250 526170 345306 526226
rect 345374 526170 345430 526226
rect 345498 526170 345554 526226
rect 345622 526170 345678 526226
rect 345250 526046 345306 526102
rect 345374 526046 345430 526102
rect 345498 526046 345554 526102
rect 345622 526046 345678 526102
rect 345250 525922 345306 525978
rect 345374 525922 345430 525978
rect 345498 525922 345554 525978
rect 345622 525922 345678 525978
rect 345250 508294 345306 508350
rect 345374 508294 345430 508350
rect 345498 508294 345554 508350
rect 345622 508294 345678 508350
rect 345250 508170 345306 508226
rect 345374 508170 345430 508226
rect 345498 508170 345554 508226
rect 345622 508170 345678 508226
rect 345250 508046 345306 508102
rect 345374 508046 345430 508102
rect 345498 508046 345554 508102
rect 345622 508046 345678 508102
rect 345250 507922 345306 507978
rect 345374 507922 345430 507978
rect 345498 507922 345554 507978
rect 345622 507922 345678 507978
rect 345250 490294 345306 490350
rect 345374 490294 345430 490350
rect 345498 490294 345554 490350
rect 345622 490294 345678 490350
rect 345250 490170 345306 490226
rect 345374 490170 345430 490226
rect 345498 490170 345554 490226
rect 345622 490170 345678 490226
rect 345250 490046 345306 490102
rect 345374 490046 345430 490102
rect 345498 490046 345554 490102
rect 345622 490046 345678 490102
rect 345250 489922 345306 489978
rect 345374 489922 345430 489978
rect 345498 489922 345554 489978
rect 345622 489922 345678 489978
rect 345250 472294 345306 472350
rect 345374 472294 345430 472350
rect 345498 472294 345554 472350
rect 345622 472294 345678 472350
rect 345250 472170 345306 472226
rect 345374 472170 345430 472226
rect 345498 472170 345554 472226
rect 345622 472170 345678 472226
rect 345250 472046 345306 472102
rect 345374 472046 345430 472102
rect 345498 472046 345554 472102
rect 345622 472046 345678 472102
rect 345250 471922 345306 471978
rect 345374 471922 345430 471978
rect 345498 471922 345554 471978
rect 345622 471922 345678 471978
rect 345250 454294 345306 454350
rect 345374 454294 345430 454350
rect 345498 454294 345554 454350
rect 345622 454294 345678 454350
rect 345250 454170 345306 454226
rect 345374 454170 345430 454226
rect 345498 454170 345554 454226
rect 345622 454170 345678 454226
rect 345250 454046 345306 454102
rect 345374 454046 345430 454102
rect 345498 454046 345554 454102
rect 345622 454046 345678 454102
rect 345250 453922 345306 453978
rect 345374 453922 345430 453978
rect 345498 453922 345554 453978
rect 345622 453922 345678 453978
rect 340998 436261 341054 436317
rect 341122 436261 341178 436317
rect 340998 436137 341054 436193
rect 341122 436137 341178 436193
rect 340998 436013 341054 436069
rect 341122 436013 341178 436069
rect 310278 435889 310334 435945
rect 310402 435889 310458 435945
rect 345250 436322 345306 436378
rect 345374 436322 345430 436378
rect 345498 436322 345554 436378
rect 345622 436322 345678 436378
rect 345250 436198 345306 436254
rect 345374 436198 345430 436254
rect 345498 436198 345554 436254
rect 345622 436198 345678 436254
rect 345250 436074 345306 436130
rect 345374 436074 345430 436130
rect 345498 436074 345554 436130
rect 345622 436074 345678 436130
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 348970 514294 349026 514350
rect 349094 514294 349150 514350
rect 349218 514294 349274 514350
rect 349342 514294 349398 514350
rect 348970 514170 349026 514226
rect 349094 514170 349150 514226
rect 349218 514170 349274 514226
rect 349342 514170 349398 514226
rect 348970 514046 349026 514102
rect 349094 514046 349150 514102
rect 349218 514046 349274 514102
rect 349342 514046 349398 514102
rect 348970 513922 349026 513978
rect 349094 513922 349150 513978
rect 349218 513922 349274 513978
rect 349342 513922 349398 513978
rect 348970 496294 349026 496350
rect 349094 496294 349150 496350
rect 349218 496294 349274 496350
rect 349342 496294 349398 496350
rect 348970 496170 349026 496226
rect 349094 496170 349150 496226
rect 349218 496170 349274 496226
rect 349342 496170 349398 496226
rect 348970 496046 349026 496102
rect 349094 496046 349150 496102
rect 349218 496046 349274 496102
rect 349342 496046 349398 496102
rect 348970 495922 349026 495978
rect 349094 495922 349150 495978
rect 349218 495922 349274 495978
rect 349342 495922 349398 495978
rect 348970 478294 349026 478350
rect 349094 478294 349150 478350
rect 349218 478294 349274 478350
rect 349342 478294 349398 478350
rect 348970 478170 349026 478226
rect 349094 478170 349150 478226
rect 349218 478170 349274 478226
rect 349342 478170 349398 478226
rect 348970 478046 349026 478102
rect 349094 478046 349150 478102
rect 349218 478046 349274 478102
rect 349342 478046 349398 478102
rect 348970 477922 349026 477978
rect 349094 477922 349150 477978
rect 349218 477922 349274 477978
rect 349342 477922 349398 477978
rect 348970 460294 349026 460350
rect 349094 460294 349150 460350
rect 349218 460294 349274 460350
rect 349342 460294 349398 460350
rect 348970 460170 349026 460226
rect 349094 460170 349150 460226
rect 349218 460170 349274 460226
rect 349342 460170 349398 460226
rect 348970 460046 349026 460102
rect 349094 460046 349150 460102
rect 349218 460046 349274 460102
rect 349342 460046 349398 460102
rect 348970 459922 349026 459978
rect 349094 459922 349150 459978
rect 349218 459922 349274 459978
rect 349342 459922 349398 459978
rect 348970 442294 349026 442350
rect 349094 442294 349150 442350
rect 349218 442294 349274 442350
rect 349342 442294 349398 442350
rect 348970 442170 349026 442226
rect 349094 442170 349150 442226
rect 349218 442170 349274 442226
rect 349342 442170 349398 442226
rect 348970 442046 349026 442102
rect 349094 442046 349150 442102
rect 349218 442046 349274 442102
rect 349342 442046 349398 442102
rect 348970 441922 349026 441978
rect 349094 441922 349150 441978
rect 349218 441922 349274 441978
rect 349342 441922 349398 441978
rect 340998 435889 341054 435945
rect 341122 435889 341178 435945
rect 79878 424294 79934 424350
rect 80002 424294 80058 424350
rect 79878 424170 79934 424226
rect 80002 424170 80058 424226
rect 79878 424046 79934 424102
rect 80002 424046 80058 424102
rect 79878 423922 79934 423978
rect 80002 423922 80058 423978
rect 110598 424294 110654 424350
rect 110722 424294 110778 424350
rect 110598 424170 110654 424226
rect 110722 424170 110778 424226
rect 110598 424046 110654 424102
rect 110722 424046 110778 424102
rect 110598 423922 110654 423978
rect 110722 423922 110778 423978
rect 141318 424294 141374 424350
rect 141442 424294 141498 424350
rect 141318 424170 141374 424226
rect 141442 424170 141498 424226
rect 141318 424046 141374 424102
rect 141442 424046 141498 424102
rect 141318 423922 141374 423978
rect 141442 423922 141498 423978
rect 172038 424294 172094 424350
rect 172162 424294 172218 424350
rect 172038 424170 172094 424226
rect 172162 424170 172218 424226
rect 172038 424046 172094 424102
rect 172162 424046 172218 424102
rect 172038 423922 172094 423978
rect 172162 423922 172218 423978
rect 202758 424294 202814 424350
rect 202882 424294 202938 424350
rect 202758 424170 202814 424226
rect 202882 424170 202938 424226
rect 202758 424046 202814 424102
rect 202882 424046 202938 424102
rect 202758 423922 202814 423978
rect 202882 423922 202938 423978
rect 233478 424294 233534 424350
rect 233602 424294 233658 424350
rect 233478 424170 233534 424226
rect 233602 424170 233658 424226
rect 233478 424046 233534 424102
rect 233602 424046 233658 424102
rect 233478 423922 233534 423978
rect 233602 423922 233658 423978
rect 264198 424294 264254 424350
rect 264322 424294 264378 424350
rect 264198 424170 264254 424226
rect 264322 424170 264378 424226
rect 264198 424046 264254 424102
rect 264322 424046 264378 424102
rect 264198 423922 264254 423978
rect 264322 423922 264378 423978
rect 294918 424294 294974 424350
rect 295042 424294 295098 424350
rect 294918 424170 294974 424226
rect 295042 424170 295098 424226
rect 294918 424046 294974 424102
rect 295042 424046 295098 424102
rect 294918 423922 294974 423978
rect 295042 423922 295098 423978
rect 325638 424294 325694 424350
rect 325762 424294 325818 424350
rect 325638 424170 325694 424226
rect 325762 424170 325818 424226
rect 325638 424046 325694 424102
rect 325762 424046 325818 424102
rect 325638 423922 325694 423978
rect 325762 423922 325818 423978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 363250 526294 363306 526350
rect 363374 526294 363430 526350
rect 363498 526294 363554 526350
rect 363622 526294 363678 526350
rect 363250 526170 363306 526226
rect 363374 526170 363430 526226
rect 363498 526170 363554 526226
rect 363622 526170 363678 526226
rect 363250 526046 363306 526102
rect 363374 526046 363430 526102
rect 363498 526046 363554 526102
rect 363622 526046 363678 526102
rect 363250 525922 363306 525978
rect 363374 525922 363430 525978
rect 363498 525922 363554 525978
rect 363622 525922 363678 525978
rect 363250 508294 363306 508350
rect 363374 508294 363430 508350
rect 363498 508294 363554 508350
rect 363622 508294 363678 508350
rect 363250 508170 363306 508226
rect 363374 508170 363430 508226
rect 363498 508170 363554 508226
rect 363622 508170 363678 508226
rect 363250 508046 363306 508102
rect 363374 508046 363430 508102
rect 363498 508046 363554 508102
rect 363622 508046 363678 508102
rect 363250 507922 363306 507978
rect 363374 507922 363430 507978
rect 363498 507922 363554 507978
rect 363622 507922 363678 507978
rect 363250 490294 363306 490350
rect 363374 490294 363430 490350
rect 363498 490294 363554 490350
rect 363622 490294 363678 490350
rect 363250 490170 363306 490226
rect 363374 490170 363430 490226
rect 363498 490170 363554 490226
rect 363622 490170 363678 490226
rect 363250 490046 363306 490102
rect 363374 490046 363430 490102
rect 363498 490046 363554 490102
rect 363622 490046 363678 490102
rect 363250 489922 363306 489978
rect 363374 489922 363430 489978
rect 363498 489922 363554 489978
rect 363622 489922 363678 489978
rect 363250 472294 363306 472350
rect 363374 472294 363430 472350
rect 363498 472294 363554 472350
rect 363622 472294 363678 472350
rect 363250 472170 363306 472226
rect 363374 472170 363430 472226
rect 363498 472170 363554 472226
rect 363622 472170 363678 472226
rect 363250 472046 363306 472102
rect 363374 472046 363430 472102
rect 363498 472046 363554 472102
rect 363622 472046 363678 472102
rect 363250 471922 363306 471978
rect 363374 471922 363430 471978
rect 363498 471922 363554 471978
rect 363622 471922 363678 471978
rect 363250 454294 363306 454350
rect 363374 454294 363430 454350
rect 363498 454294 363554 454350
rect 363622 454294 363678 454350
rect 363250 454170 363306 454226
rect 363374 454170 363430 454226
rect 363498 454170 363554 454226
rect 363622 454170 363678 454226
rect 363250 454046 363306 454102
rect 363374 454046 363430 454102
rect 363498 454046 363554 454102
rect 363622 454046 363678 454102
rect 363250 453922 363306 453978
rect 363374 453922 363430 453978
rect 363498 453922 363554 453978
rect 363622 453922 363678 453978
rect 363250 436294 363306 436350
rect 363374 436294 363430 436350
rect 363498 436294 363554 436350
rect 363622 436294 363678 436350
rect 363250 436170 363306 436226
rect 363374 436170 363430 436226
rect 363498 436170 363554 436226
rect 363622 436170 363678 436226
rect 363250 436046 363306 436102
rect 363374 436046 363430 436102
rect 363498 436046 363554 436102
rect 363622 436046 363678 436102
rect 363250 435922 363306 435978
rect 363374 435922 363430 435978
rect 363498 435922 363554 435978
rect 363622 435922 363678 435978
rect 348970 424294 349026 424350
rect 349094 424294 349150 424350
rect 349218 424294 349274 424350
rect 349342 424294 349398 424350
rect 348970 424170 349026 424226
rect 349094 424170 349150 424226
rect 349218 424170 349274 424226
rect 349342 424170 349398 424226
rect 348970 424046 349026 424102
rect 349094 424046 349150 424102
rect 349218 424046 349274 424102
rect 349342 424046 349398 424102
rect 348970 423922 349026 423978
rect 349094 423922 349150 423978
rect 349218 423922 349274 423978
rect 349342 423922 349398 423978
rect 57250 418294 57306 418350
rect 57374 418294 57430 418350
rect 57498 418294 57554 418350
rect 57622 418294 57678 418350
rect 57250 418170 57306 418226
rect 57374 418170 57430 418226
rect 57498 418170 57554 418226
rect 57622 418170 57678 418226
rect 57250 418046 57306 418102
rect 57374 418046 57430 418102
rect 57498 418046 57554 418102
rect 57622 418046 57678 418102
rect 57250 417922 57306 417978
rect 57374 417922 57430 417978
rect 57498 417922 57554 417978
rect 57622 417922 57678 417978
rect 64518 418294 64574 418350
rect 64642 418294 64698 418350
rect 64518 418170 64574 418226
rect 64642 418170 64698 418226
rect 64518 418046 64574 418102
rect 64642 418046 64698 418102
rect 64518 417922 64574 417978
rect 64642 417922 64698 417978
rect 95238 418294 95294 418350
rect 95362 418294 95418 418350
rect 95238 418170 95294 418226
rect 95362 418170 95418 418226
rect 95238 418046 95294 418102
rect 95362 418046 95418 418102
rect 95238 417922 95294 417978
rect 95362 417922 95418 417978
rect 125958 418294 126014 418350
rect 126082 418294 126138 418350
rect 125958 418170 126014 418226
rect 126082 418170 126138 418226
rect 125958 418046 126014 418102
rect 126082 418046 126138 418102
rect 125958 417922 126014 417978
rect 126082 417922 126138 417978
rect 156678 418294 156734 418350
rect 156802 418294 156858 418350
rect 156678 418170 156734 418226
rect 156802 418170 156858 418226
rect 156678 418046 156734 418102
rect 156802 418046 156858 418102
rect 156678 417922 156734 417978
rect 156802 417922 156858 417978
rect 187398 418294 187454 418350
rect 187522 418294 187578 418350
rect 187398 418170 187454 418226
rect 187522 418170 187578 418226
rect 187398 418046 187454 418102
rect 187522 418046 187578 418102
rect 187398 417922 187454 417978
rect 187522 417922 187578 417978
rect 218118 418294 218174 418350
rect 218242 418294 218298 418350
rect 218118 418170 218174 418226
rect 218242 418170 218298 418226
rect 218118 418046 218174 418102
rect 218242 418046 218298 418102
rect 218118 417922 218174 417978
rect 218242 417922 218298 417978
rect 248838 418294 248894 418350
rect 248962 418294 249018 418350
rect 248838 418170 248894 418226
rect 248962 418170 249018 418226
rect 248838 418046 248894 418102
rect 248962 418046 249018 418102
rect 248838 417922 248894 417978
rect 248962 417922 249018 417978
rect 279558 418294 279614 418350
rect 279682 418294 279738 418350
rect 279558 418170 279614 418226
rect 279682 418170 279738 418226
rect 279558 418046 279614 418102
rect 279682 418046 279738 418102
rect 279558 417922 279614 417978
rect 279682 417922 279738 417978
rect 310278 418294 310334 418350
rect 310402 418294 310458 418350
rect 310278 418170 310334 418226
rect 310402 418170 310458 418226
rect 310278 418046 310334 418102
rect 310402 418046 310458 418102
rect 310278 417922 310334 417978
rect 310402 417922 310458 417978
rect 340998 418294 341054 418350
rect 341122 418294 341178 418350
rect 340998 418170 341054 418226
rect 341122 418170 341178 418226
rect 340998 418046 341054 418102
rect 341122 418046 341178 418102
rect 340998 417922 341054 417978
rect 341122 417922 341178 417978
rect 79878 406294 79934 406350
rect 80002 406294 80058 406350
rect 79878 406170 79934 406226
rect 80002 406170 80058 406226
rect 79878 406046 79934 406102
rect 80002 406046 80058 406102
rect 79878 405922 79934 405978
rect 80002 405922 80058 405978
rect 110598 406294 110654 406350
rect 110722 406294 110778 406350
rect 110598 406170 110654 406226
rect 110722 406170 110778 406226
rect 110598 406046 110654 406102
rect 110722 406046 110778 406102
rect 110598 405922 110654 405978
rect 110722 405922 110778 405978
rect 141318 406294 141374 406350
rect 141442 406294 141498 406350
rect 141318 406170 141374 406226
rect 141442 406170 141498 406226
rect 141318 406046 141374 406102
rect 141442 406046 141498 406102
rect 141318 405922 141374 405978
rect 141442 405922 141498 405978
rect 172038 406294 172094 406350
rect 172162 406294 172218 406350
rect 172038 406170 172094 406226
rect 172162 406170 172218 406226
rect 172038 406046 172094 406102
rect 172162 406046 172218 406102
rect 172038 405922 172094 405978
rect 172162 405922 172218 405978
rect 202758 406294 202814 406350
rect 202882 406294 202938 406350
rect 202758 406170 202814 406226
rect 202882 406170 202938 406226
rect 202758 406046 202814 406102
rect 202882 406046 202938 406102
rect 202758 405922 202814 405978
rect 202882 405922 202938 405978
rect 233478 406294 233534 406350
rect 233602 406294 233658 406350
rect 233478 406170 233534 406226
rect 233602 406170 233658 406226
rect 233478 406046 233534 406102
rect 233602 406046 233658 406102
rect 233478 405922 233534 405978
rect 233602 405922 233658 405978
rect 264198 406294 264254 406350
rect 264322 406294 264378 406350
rect 264198 406170 264254 406226
rect 264322 406170 264378 406226
rect 264198 406046 264254 406102
rect 264322 406046 264378 406102
rect 264198 405922 264254 405978
rect 264322 405922 264378 405978
rect 294918 406294 294974 406350
rect 295042 406294 295098 406350
rect 294918 406170 294974 406226
rect 295042 406170 295098 406226
rect 294918 406046 294974 406102
rect 295042 406046 295098 406102
rect 294918 405922 294974 405978
rect 295042 405922 295098 405978
rect 325638 406294 325694 406350
rect 325762 406294 325818 406350
rect 325638 406170 325694 406226
rect 325762 406170 325818 406226
rect 325638 406046 325694 406102
rect 325762 406046 325818 406102
rect 325638 405922 325694 405978
rect 325762 405922 325818 405978
rect 356358 424294 356414 424350
rect 356482 424294 356538 424350
rect 356358 424170 356414 424226
rect 356482 424170 356538 424226
rect 356358 424046 356414 424102
rect 356482 424046 356538 424102
rect 356358 423922 356414 423978
rect 356482 423922 356538 423978
rect 363250 418294 363306 418350
rect 363374 418294 363430 418350
rect 363498 418294 363554 418350
rect 363622 418294 363678 418350
rect 363250 418170 363306 418226
rect 363374 418170 363430 418226
rect 363498 418170 363554 418226
rect 363622 418170 363678 418226
rect 363250 418046 363306 418102
rect 363374 418046 363430 418102
rect 363498 418046 363554 418102
rect 363622 418046 363678 418102
rect 363250 417922 363306 417978
rect 363374 417922 363430 417978
rect 363498 417922 363554 417978
rect 363622 417922 363678 417978
rect 348970 406294 349026 406350
rect 349094 406294 349150 406350
rect 349218 406294 349274 406350
rect 349342 406294 349398 406350
rect 348970 406170 349026 406226
rect 349094 406170 349150 406226
rect 349218 406170 349274 406226
rect 349342 406170 349398 406226
rect 348970 406046 349026 406102
rect 349094 406046 349150 406102
rect 349218 406046 349274 406102
rect 349342 406046 349398 406102
rect 348970 405922 349026 405978
rect 349094 405922 349150 405978
rect 349218 405922 349274 405978
rect 349342 405922 349398 405978
rect 57250 400294 57306 400350
rect 57374 400294 57430 400350
rect 57498 400294 57554 400350
rect 57622 400294 57678 400350
rect 57250 400170 57306 400226
rect 57374 400170 57430 400226
rect 57498 400170 57554 400226
rect 57622 400170 57678 400226
rect 57250 400046 57306 400102
rect 57374 400046 57430 400102
rect 57498 400046 57554 400102
rect 57622 400046 57678 400102
rect 57250 399922 57306 399978
rect 57374 399922 57430 399978
rect 57498 399922 57554 399978
rect 57622 399922 57678 399978
rect 64518 400294 64574 400350
rect 64642 400294 64698 400350
rect 64518 400170 64574 400226
rect 64642 400170 64698 400226
rect 64518 400046 64574 400102
rect 64642 400046 64698 400102
rect 64518 399922 64574 399978
rect 64642 399922 64698 399978
rect 95238 400294 95294 400350
rect 95362 400294 95418 400350
rect 95238 400170 95294 400226
rect 95362 400170 95418 400226
rect 95238 400046 95294 400102
rect 95362 400046 95418 400102
rect 95238 399922 95294 399978
rect 95362 399922 95418 399978
rect 125958 400294 126014 400350
rect 126082 400294 126138 400350
rect 125958 400170 126014 400226
rect 126082 400170 126138 400226
rect 125958 400046 126014 400102
rect 126082 400046 126138 400102
rect 125958 399922 126014 399978
rect 126082 399922 126138 399978
rect 156678 400294 156734 400350
rect 156802 400294 156858 400350
rect 156678 400170 156734 400226
rect 156802 400170 156858 400226
rect 156678 400046 156734 400102
rect 156802 400046 156858 400102
rect 156678 399922 156734 399978
rect 156802 399922 156858 399978
rect 187398 400294 187454 400350
rect 187522 400294 187578 400350
rect 187398 400170 187454 400226
rect 187522 400170 187578 400226
rect 187398 400046 187454 400102
rect 187522 400046 187578 400102
rect 187398 399922 187454 399978
rect 187522 399922 187578 399978
rect 218118 400294 218174 400350
rect 218242 400294 218298 400350
rect 218118 400170 218174 400226
rect 218242 400170 218298 400226
rect 218118 400046 218174 400102
rect 218242 400046 218298 400102
rect 218118 399922 218174 399978
rect 218242 399922 218298 399978
rect 248838 400294 248894 400350
rect 248962 400294 249018 400350
rect 248838 400170 248894 400226
rect 248962 400170 249018 400226
rect 248838 400046 248894 400102
rect 248962 400046 249018 400102
rect 248838 399922 248894 399978
rect 248962 399922 249018 399978
rect 279558 400294 279614 400350
rect 279682 400294 279738 400350
rect 279558 400170 279614 400226
rect 279682 400170 279738 400226
rect 279558 400046 279614 400102
rect 279682 400046 279738 400102
rect 279558 399922 279614 399978
rect 279682 399922 279738 399978
rect 310278 400294 310334 400350
rect 310402 400294 310458 400350
rect 310278 400170 310334 400226
rect 310402 400170 310458 400226
rect 310278 400046 310334 400102
rect 310402 400046 310458 400102
rect 310278 399922 310334 399978
rect 310402 399922 310458 399978
rect 340998 400294 341054 400350
rect 341122 400294 341178 400350
rect 340998 400170 341054 400226
rect 341122 400170 341178 400226
rect 340998 400046 341054 400102
rect 341122 400046 341178 400102
rect 340998 399922 341054 399978
rect 341122 399922 341178 399978
rect 79878 388294 79934 388350
rect 80002 388294 80058 388350
rect 79878 388170 79934 388226
rect 80002 388170 80058 388226
rect 79878 388046 79934 388102
rect 80002 388046 80058 388102
rect 79878 387922 79934 387978
rect 80002 387922 80058 387978
rect 110598 388294 110654 388350
rect 110722 388294 110778 388350
rect 110598 388170 110654 388226
rect 110722 388170 110778 388226
rect 110598 388046 110654 388102
rect 110722 388046 110778 388102
rect 110598 387922 110654 387978
rect 110722 387922 110778 387978
rect 141318 388294 141374 388350
rect 141442 388294 141498 388350
rect 141318 388170 141374 388226
rect 141442 388170 141498 388226
rect 141318 388046 141374 388102
rect 141442 388046 141498 388102
rect 141318 387922 141374 387978
rect 141442 387922 141498 387978
rect 172038 388294 172094 388350
rect 172162 388294 172218 388350
rect 172038 388170 172094 388226
rect 172162 388170 172218 388226
rect 172038 388046 172094 388102
rect 172162 388046 172218 388102
rect 172038 387922 172094 387978
rect 172162 387922 172218 387978
rect 202758 388294 202814 388350
rect 202882 388294 202938 388350
rect 202758 388170 202814 388226
rect 202882 388170 202938 388226
rect 202758 388046 202814 388102
rect 202882 388046 202938 388102
rect 202758 387922 202814 387978
rect 202882 387922 202938 387978
rect 233478 388294 233534 388350
rect 233602 388294 233658 388350
rect 233478 388170 233534 388226
rect 233602 388170 233658 388226
rect 233478 388046 233534 388102
rect 233602 388046 233658 388102
rect 233478 387922 233534 387978
rect 233602 387922 233658 387978
rect 264198 388294 264254 388350
rect 264322 388294 264378 388350
rect 264198 388170 264254 388226
rect 264322 388170 264378 388226
rect 264198 388046 264254 388102
rect 264322 388046 264378 388102
rect 264198 387922 264254 387978
rect 264322 387922 264378 387978
rect 294918 388294 294974 388350
rect 295042 388294 295098 388350
rect 294918 388170 294974 388226
rect 295042 388170 295098 388226
rect 294918 388046 294974 388102
rect 295042 388046 295098 388102
rect 294918 387922 294974 387978
rect 295042 387922 295098 387978
rect 325638 388294 325694 388350
rect 325762 388294 325818 388350
rect 325638 388170 325694 388226
rect 325762 388170 325818 388226
rect 325638 388046 325694 388102
rect 325762 388046 325818 388102
rect 325638 387922 325694 387978
rect 325762 387922 325818 387978
rect 356358 406294 356414 406350
rect 356482 406294 356538 406350
rect 356358 406170 356414 406226
rect 356482 406170 356538 406226
rect 356358 406046 356414 406102
rect 356482 406046 356538 406102
rect 356358 405922 356414 405978
rect 356482 405922 356538 405978
rect 363250 400294 363306 400350
rect 363374 400294 363430 400350
rect 363498 400294 363554 400350
rect 363622 400294 363678 400350
rect 363250 400170 363306 400226
rect 363374 400170 363430 400226
rect 363498 400170 363554 400226
rect 363622 400170 363678 400226
rect 363250 400046 363306 400102
rect 363374 400046 363430 400102
rect 363498 400046 363554 400102
rect 363622 400046 363678 400102
rect 363250 399922 363306 399978
rect 363374 399922 363430 399978
rect 363498 399922 363554 399978
rect 363622 399922 363678 399978
rect 348970 388294 349026 388350
rect 349094 388294 349150 388350
rect 349218 388294 349274 388350
rect 349342 388294 349398 388350
rect 348970 388170 349026 388226
rect 349094 388170 349150 388226
rect 349218 388170 349274 388226
rect 349342 388170 349398 388226
rect 348970 388046 349026 388102
rect 349094 388046 349150 388102
rect 349218 388046 349274 388102
rect 349342 388046 349398 388102
rect 348970 387922 349026 387978
rect 349094 387922 349150 387978
rect 349218 387922 349274 387978
rect 349342 387922 349398 387978
rect 57250 382294 57306 382350
rect 57374 382294 57430 382350
rect 57498 382294 57554 382350
rect 57622 382294 57678 382350
rect 57250 382170 57306 382226
rect 57374 382170 57430 382226
rect 57498 382170 57554 382226
rect 57622 382170 57678 382226
rect 57250 382046 57306 382102
rect 57374 382046 57430 382102
rect 57498 382046 57554 382102
rect 57622 382046 57678 382102
rect 57250 381922 57306 381978
rect 57374 381922 57430 381978
rect 57498 381922 57554 381978
rect 57622 381922 57678 381978
rect 64518 382294 64574 382350
rect 64642 382294 64698 382350
rect 64518 382170 64574 382226
rect 64642 382170 64698 382226
rect 64518 382046 64574 382102
rect 64642 382046 64698 382102
rect 64518 381922 64574 381978
rect 64642 381922 64698 381978
rect 95238 382294 95294 382350
rect 95362 382294 95418 382350
rect 95238 382170 95294 382226
rect 95362 382170 95418 382226
rect 95238 382046 95294 382102
rect 95362 382046 95418 382102
rect 95238 381922 95294 381978
rect 95362 381922 95418 381978
rect 125958 382294 126014 382350
rect 126082 382294 126138 382350
rect 125958 382170 126014 382226
rect 126082 382170 126138 382226
rect 125958 382046 126014 382102
rect 126082 382046 126138 382102
rect 125958 381922 126014 381978
rect 126082 381922 126138 381978
rect 156678 382294 156734 382350
rect 156802 382294 156858 382350
rect 156678 382170 156734 382226
rect 156802 382170 156858 382226
rect 156678 382046 156734 382102
rect 156802 382046 156858 382102
rect 156678 381922 156734 381978
rect 156802 381922 156858 381978
rect 187398 382294 187454 382350
rect 187522 382294 187578 382350
rect 187398 382170 187454 382226
rect 187522 382170 187578 382226
rect 187398 382046 187454 382102
rect 187522 382046 187578 382102
rect 187398 381922 187454 381978
rect 187522 381922 187578 381978
rect 218118 382294 218174 382350
rect 218242 382294 218298 382350
rect 218118 382170 218174 382226
rect 218242 382170 218298 382226
rect 218118 382046 218174 382102
rect 218242 382046 218298 382102
rect 218118 381922 218174 381978
rect 218242 381922 218298 381978
rect 248838 382294 248894 382350
rect 248962 382294 249018 382350
rect 248838 382170 248894 382226
rect 248962 382170 249018 382226
rect 248838 382046 248894 382102
rect 248962 382046 249018 382102
rect 248838 381922 248894 381978
rect 248962 381922 249018 381978
rect 279558 382294 279614 382350
rect 279682 382294 279738 382350
rect 279558 382170 279614 382226
rect 279682 382170 279738 382226
rect 279558 382046 279614 382102
rect 279682 382046 279738 382102
rect 279558 381922 279614 381978
rect 279682 381922 279738 381978
rect 310278 382294 310334 382350
rect 310402 382294 310458 382350
rect 310278 382170 310334 382226
rect 310402 382170 310458 382226
rect 310278 382046 310334 382102
rect 310402 382046 310458 382102
rect 310278 381922 310334 381978
rect 310402 381922 310458 381978
rect 340998 382294 341054 382350
rect 341122 382294 341178 382350
rect 340998 382170 341054 382226
rect 341122 382170 341178 382226
rect 340998 382046 341054 382102
rect 341122 382046 341178 382102
rect 340998 381922 341054 381978
rect 341122 381922 341178 381978
rect 79878 370294 79934 370350
rect 80002 370294 80058 370350
rect 79878 370170 79934 370226
rect 80002 370170 80058 370226
rect 79878 370046 79934 370102
rect 80002 370046 80058 370102
rect 79878 369922 79934 369978
rect 80002 369922 80058 369978
rect 110598 370294 110654 370350
rect 110722 370294 110778 370350
rect 110598 370170 110654 370226
rect 110722 370170 110778 370226
rect 110598 370046 110654 370102
rect 110722 370046 110778 370102
rect 110598 369922 110654 369978
rect 110722 369922 110778 369978
rect 141318 370294 141374 370350
rect 141442 370294 141498 370350
rect 141318 370170 141374 370226
rect 141442 370170 141498 370226
rect 141318 370046 141374 370102
rect 141442 370046 141498 370102
rect 141318 369922 141374 369978
rect 141442 369922 141498 369978
rect 172038 370294 172094 370350
rect 172162 370294 172218 370350
rect 172038 370170 172094 370226
rect 172162 370170 172218 370226
rect 172038 370046 172094 370102
rect 172162 370046 172218 370102
rect 172038 369922 172094 369978
rect 172162 369922 172218 369978
rect 202758 370294 202814 370350
rect 202882 370294 202938 370350
rect 202758 370170 202814 370226
rect 202882 370170 202938 370226
rect 202758 370046 202814 370102
rect 202882 370046 202938 370102
rect 202758 369922 202814 369978
rect 202882 369922 202938 369978
rect 233478 370294 233534 370350
rect 233602 370294 233658 370350
rect 233478 370170 233534 370226
rect 233602 370170 233658 370226
rect 233478 370046 233534 370102
rect 233602 370046 233658 370102
rect 233478 369922 233534 369978
rect 233602 369922 233658 369978
rect 264198 370294 264254 370350
rect 264322 370294 264378 370350
rect 264198 370170 264254 370226
rect 264322 370170 264378 370226
rect 264198 370046 264254 370102
rect 264322 370046 264378 370102
rect 264198 369922 264254 369978
rect 264322 369922 264378 369978
rect 294918 370294 294974 370350
rect 295042 370294 295098 370350
rect 294918 370170 294974 370226
rect 295042 370170 295098 370226
rect 294918 370046 294974 370102
rect 295042 370046 295098 370102
rect 294918 369922 294974 369978
rect 295042 369922 295098 369978
rect 325638 370294 325694 370350
rect 325762 370294 325818 370350
rect 325638 370170 325694 370226
rect 325762 370170 325818 370226
rect 325638 370046 325694 370102
rect 325762 370046 325818 370102
rect 325638 369922 325694 369978
rect 325762 369922 325818 369978
rect 356358 388294 356414 388350
rect 356482 388294 356538 388350
rect 356358 388170 356414 388226
rect 356482 388170 356538 388226
rect 356358 388046 356414 388102
rect 356482 388046 356538 388102
rect 356358 387922 356414 387978
rect 356482 387922 356538 387978
rect 363250 382294 363306 382350
rect 363374 382294 363430 382350
rect 363498 382294 363554 382350
rect 363622 382294 363678 382350
rect 363250 382170 363306 382226
rect 363374 382170 363430 382226
rect 363498 382170 363554 382226
rect 363622 382170 363678 382226
rect 363250 382046 363306 382102
rect 363374 382046 363430 382102
rect 363498 382046 363554 382102
rect 363622 382046 363678 382102
rect 363250 381922 363306 381978
rect 363374 381922 363430 381978
rect 363498 381922 363554 381978
rect 363622 381922 363678 381978
rect 348970 370294 349026 370350
rect 349094 370294 349150 370350
rect 349218 370294 349274 370350
rect 349342 370294 349398 370350
rect 348970 370170 349026 370226
rect 349094 370170 349150 370226
rect 349218 370170 349274 370226
rect 349342 370170 349398 370226
rect 348970 370046 349026 370102
rect 349094 370046 349150 370102
rect 349218 370046 349274 370102
rect 349342 370046 349398 370102
rect 348970 369922 349026 369978
rect 349094 369922 349150 369978
rect 349218 369922 349274 369978
rect 349342 369922 349398 369978
rect 57250 364294 57306 364350
rect 57374 364294 57430 364350
rect 57498 364294 57554 364350
rect 57622 364294 57678 364350
rect 57250 364170 57306 364226
rect 57374 364170 57430 364226
rect 57498 364170 57554 364226
rect 57622 364170 57678 364226
rect 57250 364046 57306 364102
rect 57374 364046 57430 364102
rect 57498 364046 57554 364102
rect 57622 364046 57678 364102
rect 57250 363922 57306 363978
rect 57374 363922 57430 363978
rect 57498 363922 57554 363978
rect 57622 363922 57678 363978
rect 64518 364294 64574 364350
rect 64642 364294 64698 364350
rect 64518 364170 64574 364226
rect 64642 364170 64698 364226
rect 64518 364046 64574 364102
rect 64642 364046 64698 364102
rect 64518 363922 64574 363978
rect 64642 363922 64698 363978
rect 95238 364294 95294 364350
rect 95362 364294 95418 364350
rect 95238 364170 95294 364226
rect 95362 364170 95418 364226
rect 95238 364046 95294 364102
rect 95362 364046 95418 364102
rect 95238 363922 95294 363978
rect 95362 363922 95418 363978
rect 125958 364294 126014 364350
rect 126082 364294 126138 364350
rect 125958 364170 126014 364226
rect 126082 364170 126138 364226
rect 125958 364046 126014 364102
rect 126082 364046 126138 364102
rect 125958 363922 126014 363978
rect 126082 363922 126138 363978
rect 156678 364294 156734 364350
rect 156802 364294 156858 364350
rect 156678 364170 156734 364226
rect 156802 364170 156858 364226
rect 156678 364046 156734 364102
rect 156802 364046 156858 364102
rect 156678 363922 156734 363978
rect 156802 363922 156858 363978
rect 187398 364294 187454 364350
rect 187522 364294 187578 364350
rect 187398 364170 187454 364226
rect 187522 364170 187578 364226
rect 187398 364046 187454 364102
rect 187522 364046 187578 364102
rect 187398 363922 187454 363978
rect 187522 363922 187578 363978
rect 218118 364294 218174 364350
rect 218242 364294 218298 364350
rect 218118 364170 218174 364226
rect 218242 364170 218298 364226
rect 218118 364046 218174 364102
rect 218242 364046 218298 364102
rect 218118 363922 218174 363978
rect 218242 363922 218298 363978
rect 248838 364294 248894 364350
rect 248962 364294 249018 364350
rect 248838 364170 248894 364226
rect 248962 364170 249018 364226
rect 248838 364046 248894 364102
rect 248962 364046 249018 364102
rect 248838 363922 248894 363978
rect 248962 363922 249018 363978
rect 279558 364294 279614 364350
rect 279682 364294 279738 364350
rect 279558 364170 279614 364226
rect 279682 364170 279738 364226
rect 279558 364046 279614 364102
rect 279682 364046 279738 364102
rect 279558 363922 279614 363978
rect 279682 363922 279738 363978
rect 310278 364294 310334 364350
rect 310402 364294 310458 364350
rect 310278 364170 310334 364226
rect 310402 364170 310458 364226
rect 310278 364046 310334 364102
rect 310402 364046 310458 364102
rect 310278 363922 310334 363978
rect 310402 363922 310458 363978
rect 340998 364294 341054 364350
rect 341122 364294 341178 364350
rect 340998 364170 341054 364226
rect 341122 364170 341178 364226
rect 340998 364046 341054 364102
rect 341122 364046 341178 364102
rect 340998 363922 341054 363978
rect 341122 363922 341178 363978
rect 79878 352294 79934 352350
rect 80002 352294 80058 352350
rect 79878 352170 79934 352226
rect 80002 352170 80058 352226
rect 79878 352046 79934 352102
rect 80002 352046 80058 352102
rect 79878 351922 79934 351978
rect 80002 351922 80058 351978
rect 110598 352294 110654 352350
rect 110722 352294 110778 352350
rect 110598 352170 110654 352226
rect 110722 352170 110778 352226
rect 110598 352046 110654 352102
rect 110722 352046 110778 352102
rect 110598 351922 110654 351978
rect 110722 351922 110778 351978
rect 141318 352294 141374 352350
rect 141442 352294 141498 352350
rect 141318 352170 141374 352226
rect 141442 352170 141498 352226
rect 141318 352046 141374 352102
rect 141442 352046 141498 352102
rect 141318 351922 141374 351978
rect 141442 351922 141498 351978
rect 172038 352294 172094 352350
rect 172162 352294 172218 352350
rect 172038 352170 172094 352226
rect 172162 352170 172218 352226
rect 172038 352046 172094 352102
rect 172162 352046 172218 352102
rect 172038 351922 172094 351978
rect 172162 351922 172218 351978
rect 202758 352294 202814 352350
rect 202882 352294 202938 352350
rect 202758 352170 202814 352226
rect 202882 352170 202938 352226
rect 202758 352046 202814 352102
rect 202882 352046 202938 352102
rect 202758 351922 202814 351978
rect 202882 351922 202938 351978
rect 233478 352294 233534 352350
rect 233602 352294 233658 352350
rect 233478 352170 233534 352226
rect 233602 352170 233658 352226
rect 233478 352046 233534 352102
rect 233602 352046 233658 352102
rect 233478 351922 233534 351978
rect 233602 351922 233658 351978
rect 264198 352294 264254 352350
rect 264322 352294 264378 352350
rect 264198 352170 264254 352226
rect 264322 352170 264378 352226
rect 264198 352046 264254 352102
rect 264322 352046 264378 352102
rect 264198 351922 264254 351978
rect 264322 351922 264378 351978
rect 294918 352294 294974 352350
rect 295042 352294 295098 352350
rect 294918 352170 294974 352226
rect 295042 352170 295098 352226
rect 294918 352046 294974 352102
rect 295042 352046 295098 352102
rect 294918 351922 294974 351978
rect 295042 351922 295098 351978
rect 325638 352294 325694 352350
rect 325762 352294 325818 352350
rect 325638 352170 325694 352226
rect 325762 352170 325818 352226
rect 325638 352046 325694 352102
rect 325762 352046 325818 352102
rect 325638 351922 325694 351978
rect 325762 351922 325818 351978
rect 356358 370294 356414 370350
rect 356482 370294 356538 370350
rect 356358 370170 356414 370226
rect 356482 370170 356538 370226
rect 356358 370046 356414 370102
rect 356482 370046 356538 370102
rect 356358 369922 356414 369978
rect 356482 369922 356538 369978
rect 363250 364294 363306 364350
rect 363374 364294 363430 364350
rect 363498 364294 363554 364350
rect 363622 364294 363678 364350
rect 363250 364170 363306 364226
rect 363374 364170 363430 364226
rect 363498 364170 363554 364226
rect 363622 364170 363678 364226
rect 363250 364046 363306 364102
rect 363374 364046 363430 364102
rect 363498 364046 363554 364102
rect 363622 364046 363678 364102
rect 363250 363922 363306 363978
rect 363374 363922 363430 363978
rect 363498 363922 363554 363978
rect 363622 363922 363678 363978
rect 348970 352294 349026 352350
rect 349094 352294 349150 352350
rect 349218 352294 349274 352350
rect 349342 352294 349398 352350
rect 348970 352170 349026 352226
rect 349094 352170 349150 352226
rect 349218 352170 349274 352226
rect 349342 352170 349398 352226
rect 348970 352046 349026 352102
rect 349094 352046 349150 352102
rect 349218 352046 349274 352102
rect 349342 352046 349398 352102
rect 348970 351922 349026 351978
rect 349094 351922 349150 351978
rect 349218 351922 349274 351978
rect 349342 351922 349398 351978
rect 57250 346294 57306 346350
rect 57374 346294 57430 346350
rect 57498 346294 57554 346350
rect 57622 346294 57678 346350
rect 57250 346170 57306 346226
rect 57374 346170 57430 346226
rect 57498 346170 57554 346226
rect 57622 346170 57678 346226
rect 57250 346046 57306 346102
rect 57374 346046 57430 346102
rect 57498 346046 57554 346102
rect 57622 346046 57678 346102
rect 57250 345922 57306 345978
rect 57374 345922 57430 345978
rect 57498 345922 57554 345978
rect 57622 345922 57678 345978
rect 64518 346294 64574 346350
rect 64642 346294 64698 346350
rect 64518 346170 64574 346226
rect 64642 346170 64698 346226
rect 64518 346046 64574 346102
rect 64642 346046 64698 346102
rect 64518 345922 64574 345978
rect 64642 345922 64698 345978
rect 95238 346294 95294 346350
rect 95362 346294 95418 346350
rect 95238 346170 95294 346226
rect 95362 346170 95418 346226
rect 95238 346046 95294 346102
rect 95362 346046 95418 346102
rect 95238 345922 95294 345978
rect 95362 345922 95418 345978
rect 125958 346294 126014 346350
rect 126082 346294 126138 346350
rect 125958 346170 126014 346226
rect 126082 346170 126138 346226
rect 125958 346046 126014 346102
rect 126082 346046 126138 346102
rect 125958 345922 126014 345978
rect 126082 345922 126138 345978
rect 156678 346294 156734 346350
rect 156802 346294 156858 346350
rect 156678 346170 156734 346226
rect 156802 346170 156858 346226
rect 156678 346046 156734 346102
rect 156802 346046 156858 346102
rect 156678 345922 156734 345978
rect 156802 345922 156858 345978
rect 187398 346294 187454 346350
rect 187522 346294 187578 346350
rect 187398 346170 187454 346226
rect 187522 346170 187578 346226
rect 187398 346046 187454 346102
rect 187522 346046 187578 346102
rect 187398 345922 187454 345978
rect 187522 345922 187578 345978
rect 218118 346294 218174 346350
rect 218242 346294 218298 346350
rect 218118 346170 218174 346226
rect 218242 346170 218298 346226
rect 218118 346046 218174 346102
rect 218242 346046 218298 346102
rect 218118 345922 218174 345978
rect 218242 345922 218298 345978
rect 248838 346294 248894 346350
rect 248962 346294 249018 346350
rect 248838 346170 248894 346226
rect 248962 346170 249018 346226
rect 248838 346046 248894 346102
rect 248962 346046 249018 346102
rect 248838 345922 248894 345978
rect 248962 345922 249018 345978
rect 279558 346294 279614 346350
rect 279682 346294 279738 346350
rect 279558 346170 279614 346226
rect 279682 346170 279738 346226
rect 279558 346046 279614 346102
rect 279682 346046 279738 346102
rect 279558 345922 279614 345978
rect 279682 345922 279738 345978
rect 310278 346294 310334 346350
rect 310402 346294 310458 346350
rect 310278 346170 310334 346226
rect 310402 346170 310458 346226
rect 310278 346046 310334 346102
rect 310402 346046 310458 346102
rect 310278 345922 310334 345978
rect 310402 345922 310458 345978
rect 340998 346294 341054 346350
rect 341122 346294 341178 346350
rect 340998 346170 341054 346226
rect 341122 346170 341178 346226
rect 340998 346046 341054 346102
rect 341122 346046 341178 346102
rect 340998 345922 341054 345978
rect 341122 345922 341178 345978
rect 79878 334294 79934 334350
rect 80002 334294 80058 334350
rect 79878 334170 79934 334226
rect 80002 334170 80058 334226
rect 79878 334046 79934 334102
rect 80002 334046 80058 334102
rect 79878 333922 79934 333978
rect 80002 333922 80058 333978
rect 110598 334294 110654 334350
rect 110722 334294 110778 334350
rect 110598 334170 110654 334226
rect 110722 334170 110778 334226
rect 110598 334046 110654 334102
rect 110722 334046 110778 334102
rect 110598 333922 110654 333978
rect 110722 333922 110778 333978
rect 141318 334294 141374 334350
rect 141442 334294 141498 334350
rect 141318 334170 141374 334226
rect 141442 334170 141498 334226
rect 141318 334046 141374 334102
rect 141442 334046 141498 334102
rect 141318 333922 141374 333978
rect 141442 333922 141498 333978
rect 172038 334294 172094 334350
rect 172162 334294 172218 334350
rect 172038 334170 172094 334226
rect 172162 334170 172218 334226
rect 172038 334046 172094 334102
rect 172162 334046 172218 334102
rect 172038 333922 172094 333978
rect 172162 333922 172218 333978
rect 202758 334294 202814 334350
rect 202882 334294 202938 334350
rect 202758 334170 202814 334226
rect 202882 334170 202938 334226
rect 202758 334046 202814 334102
rect 202882 334046 202938 334102
rect 202758 333922 202814 333978
rect 202882 333922 202938 333978
rect 233478 334294 233534 334350
rect 233602 334294 233658 334350
rect 233478 334170 233534 334226
rect 233602 334170 233658 334226
rect 233478 334046 233534 334102
rect 233602 334046 233658 334102
rect 233478 333922 233534 333978
rect 233602 333922 233658 333978
rect 264198 334294 264254 334350
rect 264322 334294 264378 334350
rect 264198 334170 264254 334226
rect 264322 334170 264378 334226
rect 264198 334046 264254 334102
rect 264322 334046 264378 334102
rect 264198 333922 264254 333978
rect 264322 333922 264378 333978
rect 294918 334294 294974 334350
rect 295042 334294 295098 334350
rect 294918 334170 294974 334226
rect 295042 334170 295098 334226
rect 294918 334046 294974 334102
rect 295042 334046 295098 334102
rect 294918 333922 294974 333978
rect 295042 333922 295098 333978
rect 325638 334294 325694 334350
rect 325762 334294 325818 334350
rect 325638 334170 325694 334226
rect 325762 334170 325818 334226
rect 325638 334046 325694 334102
rect 325762 334046 325818 334102
rect 325638 333922 325694 333978
rect 325762 333922 325818 333978
rect 356358 352294 356414 352350
rect 356482 352294 356538 352350
rect 356358 352170 356414 352226
rect 356482 352170 356538 352226
rect 356358 352046 356414 352102
rect 356482 352046 356538 352102
rect 356358 351922 356414 351978
rect 356482 351922 356538 351978
rect 363250 346294 363306 346350
rect 363374 346294 363430 346350
rect 363498 346294 363554 346350
rect 363622 346294 363678 346350
rect 363250 346170 363306 346226
rect 363374 346170 363430 346226
rect 363498 346170 363554 346226
rect 363622 346170 363678 346226
rect 363250 346046 363306 346102
rect 363374 346046 363430 346102
rect 363498 346046 363554 346102
rect 363622 346046 363678 346102
rect 363250 345922 363306 345978
rect 363374 345922 363430 345978
rect 363498 345922 363554 345978
rect 363622 345922 363678 345978
rect 348970 334294 349026 334350
rect 349094 334294 349150 334350
rect 349218 334294 349274 334350
rect 349342 334294 349398 334350
rect 348970 334170 349026 334226
rect 349094 334170 349150 334226
rect 349218 334170 349274 334226
rect 349342 334170 349398 334226
rect 348970 334046 349026 334102
rect 349094 334046 349150 334102
rect 349218 334046 349274 334102
rect 349342 334046 349398 334102
rect 348970 333922 349026 333978
rect 349094 333922 349150 333978
rect 349218 333922 349274 333978
rect 349342 333922 349398 333978
rect 57250 328294 57306 328350
rect 57374 328294 57430 328350
rect 57498 328294 57554 328350
rect 57622 328294 57678 328350
rect 57250 328170 57306 328226
rect 57374 328170 57430 328226
rect 57498 328170 57554 328226
rect 57622 328170 57678 328226
rect 57250 328046 57306 328102
rect 57374 328046 57430 328102
rect 57498 328046 57554 328102
rect 57622 328046 57678 328102
rect 57250 327922 57306 327978
rect 57374 327922 57430 327978
rect 57498 327922 57554 327978
rect 57622 327922 57678 327978
rect 64518 328294 64574 328350
rect 64642 328294 64698 328350
rect 64518 328170 64574 328226
rect 64642 328170 64698 328226
rect 64518 328046 64574 328102
rect 64642 328046 64698 328102
rect 64518 327922 64574 327978
rect 64642 327922 64698 327978
rect 95238 328294 95294 328350
rect 95362 328294 95418 328350
rect 95238 328170 95294 328226
rect 95362 328170 95418 328226
rect 95238 328046 95294 328102
rect 95362 328046 95418 328102
rect 95238 327922 95294 327978
rect 95362 327922 95418 327978
rect 125958 328294 126014 328350
rect 126082 328294 126138 328350
rect 125958 328170 126014 328226
rect 126082 328170 126138 328226
rect 125958 328046 126014 328102
rect 126082 328046 126138 328102
rect 125958 327922 126014 327978
rect 126082 327922 126138 327978
rect 156678 328294 156734 328350
rect 156802 328294 156858 328350
rect 156678 328170 156734 328226
rect 156802 328170 156858 328226
rect 156678 328046 156734 328102
rect 156802 328046 156858 328102
rect 156678 327922 156734 327978
rect 156802 327922 156858 327978
rect 187398 328294 187454 328350
rect 187522 328294 187578 328350
rect 187398 328170 187454 328226
rect 187522 328170 187578 328226
rect 187398 328046 187454 328102
rect 187522 328046 187578 328102
rect 187398 327922 187454 327978
rect 187522 327922 187578 327978
rect 218118 328294 218174 328350
rect 218242 328294 218298 328350
rect 218118 328170 218174 328226
rect 218242 328170 218298 328226
rect 218118 328046 218174 328102
rect 218242 328046 218298 328102
rect 218118 327922 218174 327978
rect 218242 327922 218298 327978
rect 248838 328294 248894 328350
rect 248962 328294 249018 328350
rect 248838 328170 248894 328226
rect 248962 328170 249018 328226
rect 248838 328046 248894 328102
rect 248962 328046 249018 328102
rect 248838 327922 248894 327978
rect 248962 327922 249018 327978
rect 279558 328294 279614 328350
rect 279682 328294 279738 328350
rect 279558 328170 279614 328226
rect 279682 328170 279738 328226
rect 279558 328046 279614 328102
rect 279682 328046 279738 328102
rect 279558 327922 279614 327978
rect 279682 327922 279738 327978
rect 310278 328294 310334 328350
rect 310402 328294 310458 328350
rect 310278 328170 310334 328226
rect 310402 328170 310458 328226
rect 310278 328046 310334 328102
rect 310402 328046 310458 328102
rect 310278 327922 310334 327978
rect 310402 327922 310458 327978
rect 340998 328294 341054 328350
rect 341122 328294 341178 328350
rect 340998 328170 341054 328226
rect 341122 328170 341178 328226
rect 340998 328046 341054 328102
rect 341122 328046 341178 328102
rect 340998 327922 341054 327978
rect 341122 327922 341178 327978
rect 79878 316294 79934 316350
rect 80002 316294 80058 316350
rect 79878 316170 79934 316226
rect 80002 316170 80058 316226
rect 79878 316046 79934 316102
rect 80002 316046 80058 316102
rect 79878 315922 79934 315978
rect 80002 315922 80058 315978
rect 110598 316294 110654 316350
rect 110722 316294 110778 316350
rect 110598 316170 110654 316226
rect 110722 316170 110778 316226
rect 110598 316046 110654 316102
rect 110722 316046 110778 316102
rect 110598 315922 110654 315978
rect 110722 315922 110778 315978
rect 141318 316294 141374 316350
rect 141442 316294 141498 316350
rect 141318 316170 141374 316226
rect 141442 316170 141498 316226
rect 141318 316046 141374 316102
rect 141442 316046 141498 316102
rect 141318 315922 141374 315978
rect 141442 315922 141498 315978
rect 172038 316294 172094 316350
rect 172162 316294 172218 316350
rect 172038 316170 172094 316226
rect 172162 316170 172218 316226
rect 172038 316046 172094 316102
rect 172162 316046 172218 316102
rect 172038 315922 172094 315978
rect 172162 315922 172218 315978
rect 202758 316294 202814 316350
rect 202882 316294 202938 316350
rect 202758 316170 202814 316226
rect 202882 316170 202938 316226
rect 202758 316046 202814 316102
rect 202882 316046 202938 316102
rect 202758 315922 202814 315978
rect 202882 315922 202938 315978
rect 233478 316294 233534 316350
rect 233602 316294 233658 316350
rect 233478 316170 233534 316226
rect 233602 316170 233658 316226
rect 233478 316046 233534 316102
rect 233602 316046 233658 316102
rect 233478 315922 233534 315978
rect 233602 315922 233658 315978
rect 264198 316294 264254 316350
rect 264322 316294 264378 316350
rect 264198 316170 264254 316226
rect 264322 316170 264378 316226
rect 264198 316046 264254 316102
rect 264322 316046 264378 316102
rect 264198 315922 264254 315978
rect 264322 315922 264378 315978
rect 294918 316294 294974 316350
rect 295042 316294 295098 316350
rect 294918 316170 294974 316226
rect 295042 316170 295098 316226
rect 294918 316046 294974 316102
rect 295042 316046 295098 316102
rect 294918 315922 294974 315978
rect 295042 315922 295098 315978
rect 325638 316294 325694 316350
rect 325762 316294 325818 316350
rect 325638 316170 325694 316226
rect 325762 316170 325818 316226
rect 325638 316046 325694 316102
rect 325762 316046 325818 316102
rect 325638 315922 325694 315978
rect 325762 315922 325818 315978
rect 356358 334294 356414 334350
rect 356482 334294 356538 334350
rect 356358 334170 356414 334226
rect 356482 334170 356538 334226
rect 356358 334046 356414 334102
rect 356482 334046 356538 334102
rect 356358 333922 356414 333978
rect 356482 333922 356538 333978
rect 363250 328294 363306 328350
rect 363374 328294 363430 328350
rect 363498 328294 363554 328350
rect 363622 328294 363678 328350
rect 363250 328170 363306 328226
rect 363374 328170 363430 328226
rect 363498 328170 363554 328226
rect 363622 328170 363678 328226
rect 363250 328046 363306 328102
rect 363374 328046 363430 328102
rect 363498 328046 363554 328102
rect 363622 328046 363678 328102
rect 363250 327922 363306 327978
rect 363374 327922 363430 327978
rect 363498 327922 363554 327978
rect 363622 327922 363678 327978
rect 348970 316294 349026 316350
rect 349094 316294 349150 316350
rect 349218 316294 349274 316350
rect 349342 316294 349398 316350
rect 348970 316170 349026 316226
rect 349094 316170 349150 316226
rect 349218 316170 349274 316226
rect 349342 316170 349398 316226
rect 348970 316046 349026 316102
rect 349094 316046 349150 316102
rect 349218 316046 349274 316102
rect 349342 316046 349398 316102
rect 348970 315922 349026 315978
rect 349094 315922 349150 315978
rect 349218 315922 349274 315978
rect 349342 315922 349398 315978
rect 57250 310294 57306 310350
rect 57374 310294 57430 310350
rect 57498 310294 57554 310350
rect 57622 310294 57678 310350
rect 57250 310170 57306 310226
rect 57374 310170 57430 310226
rect 57498 310170 57554 310226
rect 57622 310170 57678 310226
rect 57250 310046 57306 310102
rect 57374 310046 57430 310102
rect 57498 310046 57554 310102
rect 57622 310046 57678 310102
rect 57250 309922 57306 309978
rect 57374 309922 57430 309978
rect 57498 309922 57554 309978
rect 57622 309922 57678 309978
rect 64518 310294 64574 310350
rect 64642 310294 64698 310350
rect 64518 310170 64574 310226
rect 64642 310170 64698 310226
rect 64518 310046 64574 310102
rect 64642 310046 64698 310102
rect 64518 309922 64574 309978
rect 64642 309922 64698 309978
rect 95238 310294 95294 310350
rect 95362 310294 95418 310350
rect 95238 310170 95294 310226
rect 95362 310170 95418 310226
rect 95238 310046 95294 310102
rect 95362 310046 95418 310102
rect 95238 309922 95294 309978
rect 95362 309922 95418 309978
rect 125958 310294 126014 310350
rect 126082 310294 126138 310350
rect 125958 310170 126014 310226
rect 126082 310170 126138 310226
rect 125958 310046 126014 310102
rect 126082 310046 126138 310102
rect 125958 309922 126014 309978
rect 126082 309922 126138 309978
rect 156678 310294 156734 310350
rect 156802 310294 156858 310350
rect 156678 310170 156734 310226
rect 156802 310170 156858 310226
rect 156678 310046 156734 310102
rect 156802 310046 156858 310102
rect 156678 309922 156734 309978
rect 156802 309922 156858 309978
rect 187398 310294 187454 310350
rect 187522 310294 187578 310350
rect 187398 310170 187454 310226
rect 187522 310170 187578 310226
rect 187398 310046 187454 310102
rect 187522 310046 187578 310102
rect 187398 309922 187454 309978
rect 187522 309922 187578 309978
rect 218118 310294 218174 310350
rect 218242 310294 218298 310350
rect 218118 310170 218174 310226
rect 218242 310170 218298 310226
rect 218118 310046 218174 310102
rect 218242 310046 218298 310102
rect 218118 309922 218174 309978
rect 218242 309922 218298 309978
rect 248838 310294 248894 310350
rect 248962 310294 249018 310350
rect 248838 310170 248894 310226
rect 248962 310170 249018 310226
rect 248838 310046 248894 310102
rect 248962 310046 249018 310102
rect 248838 309922 248894 309978
rect 248962 309922 249018 309978
rect 279558 310294 279614 310350
rect 279682 310294 279738 310350
rect 279558 310170 279614 310226
rect 279682 310170 279738 310226
rect 279558 310046 279614 310102
rect 279682 310046 279738 310102
rect 279558 309922 279614 309978
rect 279682 309922 279738 309978
rect 310278 310294 310334 310350
rect 310402 310294 310458 310350
rect 310278 310170 310334 310226
rect 310402 310170 310458 310226
rect 310278 310046 310334 310102
rect 310402 310046 310458 310102
rect 310278 309922 310334 309978
rect 310402 309922 310458 309978
rect 340998 310294 341054 310350
rect 341122 310294 341178 310350
rect 340998 310170 341054 310226
rect 341122 310170 341178 310226
rect 340998 310046 341054 310102
rect 341122 310046 341178 310102
rect 340998 309922 341054 309978
rect 341122 309922 341178 309978
rect 79878 298294 79934 298350
rect 80002 298294 80058 298350
rect 79878 298170 79934 298226
rect 80002 298170 80058 298226
rect 79878 298046 79934 298102
rect 80002 298046 80058 298102
rect 79878 297922 79934 297978
rect 80002 297922 80058 297978
rect 110598 298294 110654 298350
rect 110722 298294 110778 298350
rect 110598 298170 110654 298226
rect 110722 298170 110778 298226
rect 110598 298046 110654 298102
rect 110722 298046 110778 298102
rect 110598 297922 110654 297978
rect 110722 297922 110778 297978
rect 141318 298294 141374 298350
rect 141442 298294 141498 298350
rect 141318 298170 141374 298226
rect 141442 298170 141498 298226
rect 141318 298046 141374 298102
rect 141442 298046 141498 298102
rect 141318 297922 141374 297978
rect 141442 297922 141498 297978
rect 172038 298294 172094 298350
rect 172162 298294 172218 298350
rect 172038 298170 172094 298226
rect 172162 298170 172218 298226
rect 172038 298046 172094 298102
rect 172162 298046 172218 298102
rect 172038 297922 172094 297978
rect 172162 297922 172218 297978
rect 202758 298294 202814 298350
rect 202882 298294 202938 298350
rect 202758 298170 202814 298226
rect 202882 298170 202938 298226
rect 202758 298046 202814 298102
rect 202882 298046 202938 298102
rect 202758 297922 202814 297978
rect 202882 297922 202938 297978
rect 233478 298294 233534 298350
rect 233602 298294 233658 298350
rect 233478 298170 233534 298226
rect 233602 298170 233658 298226
rect 233478 298046 233534 298102
rect 233602 298046 233658 298102
rect 233478 297922 233534 297978
rect 233602 297922 233658 297978
rect 264198 298294 264254 298350
rect 264322 298294 264378 298350
rect 264198 298170 264254 298226
rect 264322 298170 264378 298226
rect 264198 298046 264254 298102
rect 264322 298046 264378 298102
rect 264198 297922 264254 297978
rect 264322 297922 264378 297978
rect 294918 298294 294974 298350
rect 295042 298294 295098 298350
rect 294918 298170 294974 298226
rect 295042 298170 295098 298226
rect 294918 298046 294974 298102
rect 295042 298046 295098 298102
rect 294918 297922 294974 297978
rect 295042 297922 295098 297978
rect 325638 298294 325694 298350
rect 325762 298294 325818 298350
rect 325638 298170 325694 298226
rect 325762 298170 325818 298226
rect 325638 298046 325694 298102
rect 325762 298046 325818 298102
rect 325638 297922 325694 297978
rect 325762 297922 325818 297978
rect 356358 316294 356414 316350
rect 356482 316294 356538 316350
rect 356358 316170 356414 316226
rect 356482 316170 356538 316226
rect 356358 316046 356414 316102
rect 356482 316046 356538 316102
rect 356358 315922 356414 315978
rect 356482 315922 356538 315978
rect 363250 310294 363306 310350
rect 363374 310294 363430 310350
rect 363498 310294 363554 310350
rect 363622 310294 363678 310350
rect 363250 310170 363306 310226
rect 363374 310170 363430 310226
rect 363498 310170 363554 310226
rect 363622 310170 363678 310226
rect 363250 310046 363306 310102
rect 363374 310046 363430 310102
rect 363498 310046 363554 310102
rect 363622 310046 363678 310102
rect 363250 309922 363306 309978
rect 363374 309922 363430 309978
rect 363498 309922 363554 309978
rect 363622 309922 363678 309978
rect 348970 298294 349026 298350
rect 349094 298294 349150 298350
rect 349218 298294 349274 298350
rect 349342 298294 349398 298350
rect 348970 298170 349026 298226
rect 349094 298170 349150 298226
rect 349218 298170 349274 298226
rect 349342 298170 349398 298226
rect 348970 298046 349026 298102
rect 349094 298046 349150 298102
rect 349218 298046 349274 298102
rect 349342 298046 349398 298102
rect 348970 297922 349026 297978
rect 349094 297922 349150 297978
rect 349218 297922 349274 297978
rect 349342 297922 349398 297978
rect 57250 292294 57306 292350
rect 57374 292294 57430 292350
rect 57498 292294 57554 292350
rect 57622 292294 57678 292350
rect 57250 292170 57306 292226
rect 57374 292170 57430 292226
rect 57498 292170 57554 292226
rect 57622 292170 57678 292226
rect 57250 292046 57306 292102
rect 57374 292046 57430 292102
rect 57498 292046 57554 292102
rect 57622 292046 57678 292102
rect 57250 291922 57306 291978
rect 57374 291922 57430 291978
rect 57498 291922 57554 291978
rect 57622 291922 57678 291978
rect 64518 292294 64574 292350
rect 64642 292294 64698 292350
rect 64518 292170 64574 292226
rect 64642 292170 64698 292226
rect 64518 292046 64574 292102
rect 64642 292046 64698 292102
rect 64518 291922 64574 291978
rect 64642 291922 64698 291978
rect 95238 292294 95294 292350
rect 95362 292294 95418 292350
rect 95238 292170 95294 292226
rect 95362 292170 95418 292226
rect 95238 292046 95294 292102
rect 95362 292046 95418 292102
rect 95238 291922 95294 291978
rect 95362 291922 95418 291978
rect 125958 292294 126014 292350
rect 126082 292294 126138 292350
rect 125958 292170 126014 292226
rect 126082 292170 126138 292226
rect 125958 292046 126014 292102
rect 126082 292046 126138 292102
rect 125958 291922 126014 291978
rect 126082 291922 126138 291978
rect 156678 292294 156734 292350
rect 156802 292294 156858 292350
rect 156678 292170 156734 292226
rect 156802 292170 156858 292226
rect 156678 292046 156734 292102
rect 156802 292046 156858 292102
rect 156678 291922 156734 291978
rect 156802 291922 156858 291978
rect 187398 292294 187454 292350
rect 187522 292294 187578 292350
rect 187398 292170 187454 292226
rect 187522 292170 187578 292226
rect 187398 292046 187454 292102
rect 187522 292046 187578 292102
rect 187398 291922 187454 291978
rect 187522 291922 187578 291978
rect 218118 292294 218174 292350
rect 218242 292294 218298 292350
rect 218118 292170 218174 292226
rect 218242 292170 218298 292226
rect 218118 292046 218174 292102
rect 218242 292046 218298 292102
rect 218118 291922 218174 291978
rect 218242 291922 218298 291978
rect 248838 292294 248894 292350
rect 248962 292294 249018 292350
rect 248838 292170 248894 292226
rect 248962 292170 249018 292226
rect 248838 292046 248894 292102
rect 248962 292046 249018 292102
rect 248838 291922 248894 291978
rect 248962 291922 249018 291978
rect 279558 292294 279614 292350
rect 279682 292294 279738 292350
rect 279558 292170 279614 292226
rect 279682 292170 279738 292226
rect 279558 292046 279614 292102
rect 279682 292046 279738 292102
rect 279558 291922 279614 291978
rect 279682 291922 279738 291978
rect 310278 292294 310334 292350
rect 310402 292294 310458 292350
rect 310278 292170 310334 292226
rect 310402 292170 310458 292226
rect 310278 292046 310334 292102
rect 310402 292046 310458 292102
rect 310278 291922 310334 291978
rect 310402 291922 310458 291978
rect 340998 292294 341054 292350
rect 341122 292294 341178 292350
rect 340998 292170 341054 292226
rect 341122 292170 341178 292226
rect 340998 292046 341054 292102
rect 341122 292046 341178 292102
rect 340998 291922 341054 291978
rect 341122 291922 341178 291978
rect 79878 280294 79934 280350
rect 80002 280294 80058 280350
rect 79878 280170 79934 280226
rect 80002 280170 80058 280226
rect 79878 280046 79934 280102
rect 80002 280046 80058 280102
rect 79878 279922 79934 279978
rect 80002 279922 80058 279978
rect 110598 280294 110654 280350
rect 110722 280294 110778 280350
rect 110598 280170 110654 280226
rect 110722 280170 110778 280226
rect 110598 280046 110654 280102
rect 110722 280046 110778 280102
rect 110598 279922 110654 279978
rect 110722 279922 110778 279978
rect 141318 280294 141374 280350
rect 141442 280294 141498 280350
rect 141318 280170 141374 280226
rect 141442 280170 141498 280226
rect 141318 280046 141374 280102
rect 141442 280046 141498 280102
rect 141318 279922 141374 279978
rect 141442 279922 141498 279978
rect 172038 280294 172094 280350
rect 172162 280294 172218 280350
rect 172038 280170 172094 280226
rect 172162 280170 172218 280226
rect 172038 280046 172094 280102
rect 172162 280046 172218 280102
rect 172038 279922 172094 279978
rect 172162 279922 172218 279978
rect 202758 280294 202814 280350
rect 202882 280294 202938 280350
rect 202758 280170 202814 280226
rect 202882 280170 202938 280226
rect 202758 280046 202814 280102
rect 202882 280046 202938 280102
rect 202758 279922 202814 279978
rect 202882 279922 202938 279978
rect 233478 280294 233534 280350
rect 233602 280294 233658 280350
rect 233478 280170 233534 280226
rect 233602 280170 233658 280226
rect 233478 280046 233534 280102
rect 233602 280046 233658 280102
rect 233478 279922 233534 279978
rect 233602 279922 233658 279978
rect 264198 280294 264254 280350
rect 264322 280294 264378 280350
rect 264198 280170 264254 280226
rect 264322 280170 264378 280226
rect 264198 280046 264254 280102
rect 264322 280046 264378 280102
rect 264198 279922 264254 279978
rect 264322 279922 264378 279978
rect 294918 280294 294974 280350
rect 295042 280294 295098 280350
rect 294918 280170 294974 280226
rect 295042 280170 295098 280226
rect 294918 280046 294974 280102
rect 295042 280046 295098 280102
rect 294918 279922 294974 279978
rect 295042 279922 295098 279978
rect 325638 280294 325694 280350
rect 325762 280294 325818 280350
rect 325638 280170 325694 280226
rect 325762 280170 325818 280226
rect 325638 280046 325694 280102
rect 325762 280046 325818 280102
rect 325638 279922 325694 279978
rect 325762 279922 325818 279978
rect 356358 298294 356414 298350
rect 356482 298294 356538 298350
rect 356358 298170 356414 298226
rect 356482 298170 356538 298226
rect 356358 298046 356414 298102
rect 356482 298046 356538 298102
rect 356358 297922 356414 297978
rect 356482 297922 356538 297978
rect 363250 292294 363306 292350
rect 363374 292294 363430 292350
rect 363498 292294 363554 292350
rect 363622 292294 363678 292350
rect 363250 292170 363306 292226
rect 363374 292170 363430 292226
rect 363498 292170 363554 292226
rect 363622 292170 363678 292226
rect 363250 292046 363306 292102
rect 363374 292046 363430 292102
rect 363498 292046 363554 292102
rect 363622 292046 363678 292102
rect 363250 291922 363306 291978
rect 363374 291922 363430 291978
rect 363498 291922 363554 291978
rect 363622 291922 363678 291978
rect 348970 280294 349026 280350
rect 349094 280294 349150 280350
rect 349218 280294 349274 280350
rect 349342 280294 349398 280350
rect 348970 280170 349026 280226
rect 349094 280170 349150 280226
rect 349218 280170 349274 280226
rect 349342 280170 349398 280226
rect 348970 280046 349026 280102
rect 349094 280046 349150 280102
rect 349218 280046 349274 280102
rect 349342 280046 349398 280102
rect 348970 279922 349026 279978
rect 349094 279922 349150 279978
rect 349218 279922 349274 279978
rect 349342 279922 349398 279978
rect 57250 274294 57306 274350
rect 57374 274294 57430 274350
rect 57498 274294 57554 274350
rect 57622 274294 57678 274350
rect 57250 274170 57306 274226
rect 57374 274170 57430 274226
rect 57498 274170 57554 274226
rect 57622 274170 57678 274226
rect 57250 274046 57306 274102
rect 57374 274046 57430 274102
rect 57498 274046 57554 274102
rect 57622 274046 57678 274102
rect 57250 273922 57306 273978
rect 57374 273922 57430 273978
rect 57498 273922 57554 273978
rect 57622 273922 57678 273978
rect 64518 274294 64574 274350
rect 64642 274294 64698 274350
rect 64518 274170 64574 274226
rect 64642 274170 64698 274226
rect 64518 274046 64574 274102
rect 64642 274046 64698 274102
rect 64518 273922 64574 273978
rect 64642 273922 64698 273978
rect 95238 274294 95294 274350
rect 95362 274294 95418 274350
rect 95238 274170 95294 274226
rect 95362 274170 95418 274226
rect 95238 274046 95294 274102
rect 95362 274046 95418 274102
rect 95238 273922 95294 273978
rect 95362 273922 95418 273978
rect 125958 274294 126014 274350
rect 126082 274294 126138 274350
rect 125958 274170 126014 274226
rect 126082 274170 126138 274226
rect 125958 274046 126014 274102
rect 126082 274046 126138 274102
rect 125958 273922 126014 273978
rect 126082 273922 126138 273978
rect 156678 274294 156734 274350
rect 156802 274294 156858 274350
rect 156678 274170 156734 274226
rect 156802 274170 156858 274226
rect 156678 274046 156734 274102
rect 156802 274046 156858 274102
rect 156678 273922 156734 273978
rect 156802 273922 156858 273978
rect 187398 274294 187454 274350
rect 187522 274294 187578 274350
rect 187398 274170 187454 274226
rect 187522 274170 187578 274226
rect 187398 274046 187454 274102
rect 187522 274046 187578 274102
rect 187398 273922 187454 273978
rect 187522 273922 187578 273978
rect 218118 274294 218174 274350
rect 218242 274294 218298 274350
rect 218118 274170 218174 274226
rect 218242 274170 218298 274226
rect 218118 274046 218174 274102
rect 218242 274046 218298 274102
rect 218118 273922 218174 273978
rect 218242 273922 218298 273978
rect 248838 274294 248894 274350
rect 248962 274294 249018 274350
rect 248838 274170 248894 274226
rect 248962 274170 249018 274226
rect 248838 274046 248894 274102
rect 248962 274046 249018 274102
rect 248838 273922 248894 273978
rect 248962 273922 249018 273978
rect 279558 274294 279614 274350
rect 279682 274294 279738 274350
rect 279558 274170 279614 274226
rect 279682 274170 279738 274226
rect 279558 274046 279614 274102
rect 279682 274046 279738 274102
rect 279558 273922 279614 273978
rect 279682 273922 279738 273978
rect 310278 274294 310334 274350
rect 310402 274294 310458 274350
rect 310278 274170 310334 274226
rect 310402 274170 310458 274226
rect 310278 274046 310334 274102
rect 310402 274046 310458 274102
rect 310278 273922 310334 273978
rect 310402 273922 310458 273978
rect 340998 274294 341054 274350
rect 341122 274294 341178 274350
rect 340998 274170 341054 274226
rect 341122 274170 341178 274226
rect 340998 274046 341054 274102
rect 341122 274046 341178 274102
rect 340998 273922 341054 273978
rect 341122 273922 341178 273978
rect 79878 262294 79934 262350
rect 80002 262294 80058 262350
rect 79878 262170 79934 262226
rect 80002 262170 80058 262226
rect 79878 262046 79934 262102
rect 80002 262046 80058 262102
rect 79878 261922 79934 261978
rect 80002 261922 80058 261978
rect 110598 262294 110654 262350
rect 110722 262294 110778 262350
rect 110598 262170 110654 262226
rect 110722 262170 110778 262226
rect 110598 262046 110654 262102
rect 110722 262046 110778 262102
rect 110598 261922 110654 261978
rect 110722 261922 110778 261978
rect 141318 262294 141374 262350
rect 141442 262294 141498 262350
rect 141318 262170 141374 262226
rect 141442 262170 141498 262226
rect 141318 262046 141374 262102
rect 141442 262046 141498 262102
rect 141318 261922 141374 261978
rect 141442 261922 141498 261978
rect 172038 262294 172094 262350
rect 172162 262294 172218 262350
rect 172038 262170 172094 262226
rect 172162 262170 172218 262226
rect 172038 262046 172094 262102
rect 172162 262046 172218 262102
rect 172038 261922 172094 261978
rect 172162 261922 172218 261978
rect 202758 262294 202814 262350
rect 202882 262294 202938 262350
rect 202758 262170 202814 262226
rect 202882 262170 202938 262226
rect 202758 262046 202814 262102
rect 202882 262046 202938 262102
rect 202758 261922 202814 261978
rect 202882 261922 202938 261978
rect 233478 262294 233534 262350
rect 233602 262294 233658 262350
rect 233478 262170 233534 262226
rect 233602 262170 233658 262226
rect 233478 262046 233534 262102
rect 233602 262046 233658 262102
rect 233478 261922 233534 261978
rect 233602 261922 233658 261978
rect 264198 262294 264254 262350
rect 264322 262294 264378 262350
rect 264198 262170 264254 262226
rect 264322 262170 264378 262226
rect 264198 262046 264254 262102
rect 264322 262046 264378 262102
rect 264198 261922 264254 261978
rect 264322 261922 264378 261978
rect 294918 262294 294974 262350
rect 295042 262294 295098 262350
rect 294918 262170 294974 262226
rect 295042 262170 295098 262226
rect 294918 262046 294974 262102
rect 295042 262046 295098 262102
rect 294918 261922 294974 261978
rect 295042 261922 295098 261978
rect 325638 262294 325694 262350
rect 325762 262294 325818 262350
rect 325638 262170 325694 262226
rect 325762 262170 325818 262226
rect 325638 262046 325694 262102
rect 325762 262046 325818 262102
rect 325638 261922 325694 261978
rect 325762 261922 325818 261978
rect 356358 280294 356414 280350
rect 356482 280294 356538 280350
rect 356358 280170 356414 280226
rect 356482 280170 356538 280226
rect 356358 280046 356414 280102
rect 356482 280046 356538 280102
rect 356358 279922 356414 279978
rect 356482 279922 356538 279978
rect 363250 274294 363306 274350
rect 363374 274294 363430 274350
rect 363498 274294 363554 274350
rect 363622 274294 363678 274350
rect 363250 274170 363306 274226
rect 363374 274170 363430 274226
rect 363498 274170 363554 274226
rect 363622 274170 363678 274226
rect 363250 274046 363306 274102
rect 363374 274046 363430 274102
rect 363498 274046 363554 274102
rect 363622 274046 363678 274102
rect 363250 273922 363306 273978
rect 363374 273922 363430 273978
rect 363498 273922 363554 273978
rect 363622 273922 363678 273978
rect 348970 262294 349026 262350
rect 349094 262294 349150 262350
rect 349218 262294 349274 262350
rect 349342 262294 349398 262350
rect 348970 262170 349026 262226
rect 349094 262170 349150 262226
rect 349218 262170 349274 262226
rect 349342 262170 349398 262226
rect 348970 262046 349026 262102
rect 349094 262046 349150 262102
rect 349218 262046 349274 262102
rect 349342 262046 349398 262102
rect 348970 261922 349026 261978
rect 349094 261922 349150 261978
rect 349218 261922 349274 261978
rect 349342 261922 349398 261978
rect 57250 256294 57306 256350
rect 57374 256294 57430 256350
rect 57498 256294 57554 256350
rect 57622 256294 57678 256350
rect 57250 256170 57306 256226
rect 57374 256170 57430 256226
rect 57498 256170 57554 256226
rect 57622 256170 57678 256226
rect 57250 256046 57306 256102
rect 57374 256046 57430 256102
rect 57498 256046 57554 256102
rect 57622 256046 57678 256102
rect 57250 255922 57306 255978
rect 57374 255922 57430 255978
rect 57498 255922 57554 255978
rect 57622 255922 57678 255978
rect 64518 256294 64574 256350
rect 64642 256294 64698 256350
rect 64518 256170 64574 256226
rect 64642 256170 64698 256226
rect 64518 256046 64574 256102
rect 64642 256046 64698 256102
rect 64518 255922 64574 255978
rect 64642 255922 64698 255978
rect 95238 256294 95294 256350
rect 95362 256294 95418 256350
rect 95238 256170 95294 256226
rect 95362 256170 95418 256226
rect 95238 256046 95294 256102
rect 95362 256046 95418 256102
rect 95238 255922 95294 255978
rect 95362 255922 95418 255978
rect 125958 256294 126014 256350
rect 126082 256294 126138 256350
rect 125958 256170 126014 256226
rect 126082 256170 126138 256226
rect 125958 256046 126014 256102
rect 126082 256046 126138 256102
rect 125958 255922 126014 255978
rect 126082 255922 126138 255978
rect 156678 256294 156734 256350
rect 156802 256294 156858 256350
rect 156678 256170 156734 256226
rect 156802 256170 156858 256226
rect 156678 256046 156734 256102
rect 156802 256046 156858 256102
rect 156678 255922 156734 255978
rect 156802 255922 156858 255978
rect 187398 256294 187454 256350
rect 187522 256294 187578 256350
rect 187398 256170 187454 256226
rect 187522 256170 187578 256226
rect 187398 256046 187454 256102
rect 187522 256046 187578 256102
rect 187398 255922 187454 255978
rect 187522 255922 187578 255978
rect 218118 256294 218174 256350
rect 218242 256294 218298 256350
rect 218118 256170 218174 256226
rect 218242 256170 218298 256226
rect 218118 256046 218174 256102
rect 218242 256046 218298 256102
rect 218118 255922 218174 255978
rect 218242 255922 218298 255978
rect 248838 256294 248894 256350
rect 248962 256294 249018 256350
rect 248838 256170 248894 256226
rect 248962 256170 249018 256226
rect 248838 256046 248894 256102
rect 248962 256046 249018 256102
rect 248838 255922 248894 255978
rect 248962 255922 249018 255978
rect 279558 256294 279614 256350
rect 279682 256294 279738 256350
rect 279558 256170 279614 256226
rect 279682 256170 279738 256226
rect 279558 256046 279614 256102
rect 279682 256046 279738 256102
rect 279558 255922 279614 255978
rect 279682 255922 279738 255978
rect 310278 256294 310334 256350
rect 310402 256294 310458 256350
rect 310278 256170 310334 256226
rect 310402 256170 310458 256226
rect 310278 256046 310334 256102
rect 310402 256046 310458 256102
rect 310278 255922 310334 255978
rect 310402 255922 310458 255978
rect 340998 256294 341054 256350
rect 341122 256294 341178 256350
rect 340998 256170 341054 256226
rect 341122 256170 341178 256226
rect 340998 256046 341054 256102
rect 341122 256046 341178 256102
rect 340998 255922 341054 255978
rect 341122 255922 341178 255978
rect 79878 244294 79934 244350
rect 80002 244294 80058 244350
rect 79878 244170 79934 244226
rect 80002 244170 80058 244226
rect 79878 244046 79934 244102
rect 80002 244046 80058 244102
rect 79878 243922 79934 243978
rect 80002 243922 80058 243978
rect 110598 244294 110654 244350
rect 110722 244294 110778 244350
rect 110598 244170 110654 244226
rect 110722 244170 110778 244226
rect 110598 244046 110654 244102
rect 110722 244046 110778 244102
rect 110598 243922 110654 243978
rect 110722 243922 110778 243978
rect 141318 244294 141374 244350
rect 141442 244294 141498 244350
rect 141318 244170 141374 244226
rect 141442 244170 141498 244226
rect 141318 244046 141374 244102
rect 141442 244046 141498 244102
rect 141318 243922 141374 243978
rect 141442 243922 141498 243978
rect 172038 244294 172094 244350
rect 172162 244294 172218 244350
rect 172038 244170 172094 244226
rect 172162 244170 172218 244226
rect 172038 244046 172094 244102
rect 172162 244046 172218 244102
rect 172038 243922 172094 243978
rect 172162 243922 172218 243978
rect 202758 244294 202814 244350
rect 202882 244294 202938 244350
rect 202758 244170 202814 244226
rect 202882 244170 202938 244226
rect 202758 244046 202814 244102
rect 202882 244046 202938 244102
rect 202758 243922 202814 243978
rect 202882 243922 202938 243978
rect 233478 244294 233534 244350
rect 233602 244294 233658 244350
rect 233478 244170 233534 244226
rect 233602 244170 233658 244226
rect 233478 244046 233534 244102
rect 233602 244046 233658 244102
rect 233478 243922 233534 243978
rect 233602 243922 233658 243978
rect 264198 244294 264254 244350
rect 264322 244294 264378 244350
rect 264198 244170 264254 244226
rect 264322 244170 264378 244226
rect 264198 244046 264254 244102
rect 264322 244046 264378 244102
rect 264198 243922 264254 243978
rect 264322 243922 264378 243978
rect 294918 244294 294974 244350
rect 295042 244294 295098 244350
rect 294918 244170 294974 244226
rect 295042 244170 295098 244226
rect 294918 244046 294974 244102
rect 295042 244046 295098 244102
rect 294918 243922 294974 243978
rect 295042 243922 295098 243978
rect 325638 244294 325694 244350
rect 325762 244294 325818 244350
rect 325638 244170 325694 244226
rect 325762 244170 325818 244226
rect 325638 244046 325694 244102
rect 325762 244046 325818 244102
rect 325638 243922 325694 243978
rect 325762 243922 325818 243978
rect 356358 262294 356414 262350
rect 356482 262294 356538 262350
rect 356358 262170 356414 262226
rect 356482 262170 356538 262226
rect 356358 262046 356414 262102
rect 356482 262046 356538 262102
rect 356358 261922 356414 261978
rect 356482 261922 356538 261978
rect 363250 256294 363306 256350
rect 363374 256294 363430 256350
rect 363498 256294 363554 256350
rect 363622 256294 363678 256350
rect 363250 256170 363306 256226
rect 363374 256170 363430 256226
rect 363498 256170 363554 256226
rect 363622 256170 363678 256226
rect 363250 256046 363306 256102
rect 363374 256046 363430 256102
rect 363498 256046 363554 256102
rect 363622 256046 363678 256102
rect 363250 255922 363306 255978
rect 363374 255922 363430 255978
rect 363498 255922 363554 255978
rect 363622 255922 363678 255978
rect 348970 244294 349026 244350
rect 349094 244294 349150 244350
rect 349218 244294 349274 244350
rect 349342 244294 349398 244350
rect 348970 244170 349026 244226
rect 349094 244170 349150 244226
rect 349218 244170 349274 244226
rect 349342 244170 349398 244226
rect 348970 244046 349026 244102
rect 349094 244046 349150 244102
rect 349218 244046 349274 244102
rect 349342 244046 349398 244102
rect 348970 243922 349026 243978
rect 349094 243922 349150 243978
rect 349218 243922 349274 243978
rect 349342 243922 349398 243978
rect 57250 238294 57306 238350
rect 57374 238294 57430 238350
rect 57498 238294 57554 238350
rect 57622 238294 57678 238350
rect 57250 238170 57306 238226
rect 57374 238170 57430 238226
rect 57498 238170 57554 238226
rect 57622 238170 57678 238226
rect 57250 238046 57306 238102
rect 57374 238046 57430 238102
rect 57498 238046 57554 238102
rect 57622 238046 57678 238102
rect 57250 237922 57306 237978
rect 57374 237922 57430 237978
rect 57498 237922 57554 237978
rect 57622 237922 57678 237978
rect 64518 238294 64574 238350
rect 64642 238294 64698 238350
rect 64518 238170 64574 238226
rect 64642 238170 64698 238226
rect 64518 238046 64574 238102
rect 64642 238046 64698 238102
rect 64518 237922 64574 237978
rect 64642 237922 64698 237978
rect 95238 238294 95294 238350
rect 95362 238294 95418 238350
rect 95238 238170 95294 238226
rect 95362 238170 95418 238226
rect 95238 238046 95294 238102
rect 95362 238046 95418 238102
rect 95238 237922 95294 237978
rect 95362 237922 95418 237978
rect 125958 238294 126014 238350
rect 126082 238294 126138 238350
rect 125958 238170 126014 238226
rect 126082 238170 126138 238226
rect 125958 238046 126014 238102
rect 126082 238046 126138 238102
rect 125958 237922 126014 237978
rect 126082 237922 126138 237978
rect 156678 238294 156734 238350
rect 156802 238294 156858 238350
rect 156678 238170 156734 238226
rect 156802 238170 156858 238226
rect 156678 238046 156734 238102
rect 156802 238046 156858 238102
rect 156678 237922 156734 237978
rect 156802 237922 156858 237978
rect 187398 238294 187454 238350
rect 187522 238294 187578 238350
rect 187398 238170 187454 238226
rect 187522 238170 187578 238226
rect 187398 238046 187454 238102
rect 187522 238046 187578 238102
rect 187398 237922 187454 237978
rect 187522 237922 187578 237978
rect 218118 238294 218174 238350
rect 218242 238294 218298 238350
rect 218118 238170 218174 238226
rect 218242 238170 218298 238226
rect 218118 238046 218174 238102
rect 218242 238046 218298 238102
rect 218118 237922 218174 237978
rect 218242 237922 218298 237978
rect 248838 238294 248894 238350
rect 248962 238294 249018 238350
rect 248838 238170 248894 238226
rect 248962 238170 249018 238226
rect 248838 238046 248894 238102
rect 248962 238046 249018 238102
rect 248838 237922 248894 237978
rect 248962 237922 249018 237978
rect 279558 238294 279614 238350
rect 279682 238294 279738 238350
rect 279558 238170 279614 238226
rect 279682 238170 279738 238226
rect 279558 238046 279614 238102
rect 279682 238046 279738 238102
rect 279558 237922 279614 237978
rect 279682 237922 279738 237978
rect 310278 238294 310334 238350
rect 310402 238294 310458 238350
rect 310278 238170 310334 238226
rect 310402 238170 310458 238226
rect 310278 238046 310334 238102
rect 310402 238046 310458 238102
rect 310278 237922 310334 237978
rect 310402 237922 310458 237978
rect 340998 238294 341054 238350
rect 341122 238294 341178 238350
rect 340998 238170 341054 238226
rect 341122 238170 341178 238226
rect 340998 238046 341054 238102
rect 341122 238046 341178 238102
rect 340998 237922 341054 237978
rect 341122 237922 341178 237978
rect 79878 226294 79934 226350
rect 80002 226294 80058 226350
rect 79878 226170 79934 226226
rect 80002 226170 80058 226226
rect 79878 226046 79934 226102
rect 80002 226046 80058 226102
rect 79878 225922 79934 225978
rect 80002 225922 80058 225978
rect 110598 226294 110654 226350
rect 110722 226294 110778 226350
rect 110598 226170 110654 226226
rect 110722 226170 110778 226226
rect 110598 226046 110654 226102
rect 110722 226046 110778 226102
rect 110598 225922 110654 225978
rect 110722 225922 110778 225978
rect 141318 226294 141374 226350
rect 141442 226294 141498 226350
rect 141318 226170 141374 226226
rect 141442 226170 141498 226226
rect 141318 226046 141374 226102
rect 141442 226046 141498 226102
rect 141318 225922 141374 225978
rect 141442 225922 141498 225978
rect 172038 226294 172094 226350
rect 172162 226294 172218 226350
rect 172038 226170 172094 226226
rect 172162 226170 172218 226226
rect 172038 226046 172094 226102
rect 172162 226046 172218 226102
rect 172038 225922 172094 225978
rect 172162 225922 172218 225978
rect 202758 226294 202814 226350
rect 202882 226294 202938 226350
rect 202758 226170 202814 226226
rect 202882 226170 202938 226226
rect 202758 226046 202814 226102
rect 202882 226046 202938 226102
rect 202758 225922 202814 225978
rect 202882 225922 202938 225978
rect 233478 226294 233534 226350
rect 233602 226294 233658 226350
rect 233478 226170 233534 226226
rect 233602 226170 233658 226226
rect 233478 226046 233534 226102
rect 233602 226046 233658 226102
rect 233478 225922 233534 225978
rect 233602 225922 233658 225978
rect 264198 226294 264254 226350
rect 264322 226294 264378 226350
rect 264198 226170 264254 226226
rect 264322 226170 264378 226226
rect 264198 226046 264254 226102
rect 264322 226046 264378 226102
rect 264198 225922 264254 225978
rect 264322 225922 264378 225978
rect 294918 226294 294974 226350
rect 295042 226294 295098 226350
rect 294918 226170 294974 226226
rect 295042 226170 295098 226226
rect 294918 226046 294974 226102
rect 295042 226046 295098 226102
rect 294918 225922 294974 225978
rect 295042 225922 295098 225978
rect 325638 226294 325694 226350
rect 325762 226294 325818 226350
rect 325638 226170 325694 226226
rect 325762 226170 325818 226226
rect 325638 226046 325694 226102
rect 325762 226046 325818 226102
rect 325638 225922 325694 225978
rect 325762 225922 325818 225978
rect 356358 244294 356414 244350
rect 356482 244294 356538 244350
rect 356358 244170 356414 244226
rect 356482 244170 356538 244226
rect 356358 244046 356414 244102
rect 356482 244046 356538 244102
rect 356358 243922 356414 243978
rect 356482 243922 356538 243978
rect 363250 238294 363306 238350
rect 363374 238294 363430 238350
rect 363498 238294 363554 238350
rect 363622 238294 363678 238350
rect 363250 238170 363306 238226
rect 363374 238170 363430 238226
rect 363498 238170 363554 238226
rect 363622 238170 363678 238226
rect 363250 238046 363306 238102
rect 363374 238046 363430 238102
rect 363498 238046 363554 238102
rect 363622 238046 363678 238102
rect 363250 237922 363306 237978
rect 363374 237922 363430 237978
rect 363498 237922 363554 237978
rect 363622 237922 363678 237978
rect 348970 226294 349026 226350
rect 349094 226294 349150 226350
rect 349218 226294 349274 226350
rect 349342 226294 349398 226350
rect 348970 226170 349026 226226
rect 349094 226170 349150 226226
rect 349218 226170 349274 226226
rect 349342 226170 349398 226226
rect 348970 226046 349026 226102
rect 349094 226046 349150 226102
rect 349218 226046 349274 226102
rect 349342 226046 349398 226102
rect 348970 225922 349026 225978
rect 349094 225922 349150 225978
rect 349218 225922 349274 225978
rect 349342 225922 349398 225978
rect 57250 220294 57306 220350
rect 57374 220294 57430 220350
rect 57498 220294 57554 220350
rect 57622 220294 57678 220350
rect 57250 220170 57306 220226
rect 57374 220170 57430 220226
rect 57498 220170 57554 220226
rect 57622 220170 57678 220226
rect 57250 220046 57306 220102
rect 57374 220046 57430 220102
rect 57498 220046 57554 220102
rect 57622 220046 57678 220102
rect 57250 219922 57306 219978
rect 57374 219922 57430 219978
rect 57498 219922 57554 219978
rect 57622 219922 57678 219978
rect 64518 220294 64574 220350
rect 64642 220294 64698 220350
rect 64518 220170 64574 220226
rect 64642 220170 64698 220226
rect 64518 220046 64574 220102
rect 64642 220046 64698 220102
rect 64518 219922 64574 219978
rect 64642 219922 64698 219978
rect 95238 220294 95294 220350
rect 95362 220294 95418 220350
rect 95238 220170 95294 220226
rect 95362 220170 95418 220226
rect 95238 220046 95294 220102
rect 95362 220046 95418 220102
rect 95238 219922 95294 219978
rect 95362 219922 95418 219978
rect 125958 220294 126014 220350
rect 126082 220294 126138 220350
rect 125958 220170 126014 220226
rect 126082 220170 126138 220226
rect 125958 220046 126014 220102
rect 126082 220046 126138 220102
rect 125958 219922 126014 219978
rect 126082 219922 126138 219978
rect 156678 220294 156734 220350
rect 156802 220294 156858 220350
rect 156678 220170 156734 220226
rect 156802 220170 156858 220226
rect 156678 220046 156734 220102
rect 156802 220046 156858 220102
rect 156678 219922 156734 219978
rect 156802 219922 156858 219978
rect 187398 220294 187454 220350
rect 187522 220294 187578 220350
rect 187398 220170 187454 220226
rect 187522 220170 187578 220226
rect 187398 220046 187454 220102
rect 187522 220046 187578 220102
rect 187398 219922 187454 219978
rect 187522 219922 187578 219978
rect 218118 220294 218174 220350
rect 218242 220294 218298 220350
rect 218118 220170 218174 220226
rect 218242 220170 218298 220226
rect 218118 220046 218174 220102
rect 218242 220046 218298 220102
rect 218118 219922 218174 219978
rect 218242 219922 218298 219978
rect 248838 220294 248894 220350
rect 248962 220294 249018 220350
rect 248838 220170 248894 220226
rect 248962 220170 249018 220226
rect 248838 220046 248894 220102
rect 248962 220046 249018 220102
rect 248838 219922 248894 219978
rect 248962 219922 249018 219978
rect 279558 220294 279614 220350
rect 279682 220294 279738 220350
rect 279558 220170 279614 220226
rect 279682 220170 279738 220226
rect 279558 220046 279614 220102
rect 279682 220046 279738 220102
rect 279558 219922 279614 219978
rect 279682 219922 279738 219978
rect 310278 220294 310334 220350
rect 310402 220294 310458 220350
rect 310278 220170 310334 220226
rect 310402 220170 310458 220226
rect 310278 220046 310334 220102
rect 310402 220046 310458 220102
rect 310278 219922 310334 219978
rect 310402 219922 310458 219978
rect 340998 220294 341054 220350
rect 341122 220294 341178 220350
rect 340998 220170 341054 220226
rect 341122 220170 341178 220226
rect 340998 220046 341054 220102
rect 341122 220046 341178 220102
rect 340998 219922 341054 219978
rect 341122 219922 341178 219978
rect 79878 208294 79934 208350
rect 80002 208294 80058 208350
rect 79878 208170 79934 208226
rect 80002 208170 80058 208226
rect 79878 208046 79934 208102
rect 80002 208046 80058 208102
rect 79878 207922 79934 207978
rect 80002 207922 80058 207978
rect 110598 208294 110654 208350
rect 110722 208294 110778 208350
rect 110598 208170 110654 208226
rect 110722 208170 110778 208226
rect 110598 208046 110654 208102
rect 110722 208046 110778 208102
rect 110598 207922 110654 207978
rect 110722 207922 110778 207978
rect 141318 208294 141374 208350
rect 141442 208294 141498 208350
rect 141318 208170 141374 208226
rect 141442 208170 141498 208226
rect 141318 208046 141374 208102
rect 141442 208046 141498 208102
rect 141318 207922 141374 207978
rect 141442 207922 141498 207978
rect 172038 208294 172094 208350
rect 172162 208294 172218 208350
rect 172038 208170 172094 208226
rect 172162 208170 172218 208226
rect 172038 208046 172094 208102
rect 172162 208046 172218 208102
rect 172038 207922 172094 207978
rect 172162 207922 172218 207978
rect 202758 208294 202814 208350
rect 202882 208294 202938 208350
rect 202758 208170 202814 208226
rect 202882 208170 202938 208226
rect 202758 208046 202814 208102
rect 202882 208046 202938 208102
rect 202758 207922 202814 207978
rect 202882 207922 202938 207978
rect 233478 208294 233534 208350
rect 233602 208294 233658 208350
rect 233478 208170 233534 208226
rect 233602 208170 233658 208226
rect 233478 208046 233534 208102
rect 233602 208046 233658 208102
rect 233478 207922 233534 207978
rect 233602 207922 233658 207978
rect 264198 208294 264254 208350
rect 264322 208294 264378 208350
rect 264198 208170 264254 208226
rect 264322 208170 264378 208226
rect 264198 208046 264254 208102
rect 264322 208046 264378 208102
rect 264198 207922 264254 207978
rect 264322 207922 264378 207978
rect 294918 208294 294974 208350
rect 295042 208294 295098 208350
rect 294918 208170 294974 208226
rect 295042 208170 295098 208226
rect 294918 208046 294974 208102
rect 295042 208046 295098 208102
rect 294918 207922 294974 207978
rect 295042 207922 295098 207978
rect 325638 208294 325694 208350
rect 325762 208294 325818 208350
rect 325638 208170 325694 208226
rect 325762 208170 325818 208226
rect 325638 208046 325694 208102
rect 325762 208046 325818 208102
rect 325638 207922 325694 207978
rect 325762 207922 325818 207978
rect 356358 226294 356414 226350
rect 356482 226294 356538 226350
rect 356358 226170 356414 226226
rect 356482 226170 356538 226226
rect 356358 226046 356414 226102
rect 356482 226046 356538 226102
rect 356358 225922 356414 225978
rect 356482 225922 356538 225978
rect 363250 220294 363306 220350
rect 363374 220294 363430 220350
rect 363498 220294 363554 220350
rect 363622 220294 363678 220350
rect 363250 220170 363306 220226
rect 363374 220170 363430 220226
rect 363498 220170 363554 220226
rect 363622 220170 363678 220226
rect 363250 220046 363306 220102
rect 363374 220046 363430 220102
rect 363498 220046 363554 220102
rect 363622 220046 363678 220102
rect 363250 219922 363306 219978
rect 363374 219922 363430 219978
rect 363498 219922 363554 219978
rect 363622 219922 363678 219978
rect 348970 208294 349026 208350
rect 349094 208294 349150 208350
rect 349218 208294 349274 208350
rect 349342 208294 349398 208350
rect 348970 208170 349026 208226
rect 349094 208170 349150 208226
rect 349218 208170 349274 208226
rect 349342 208170 349398 208226
rect 348970 208046 349026 208102
rect 349094 208046 349150 208102
rect 349218 208046 349274 208102
rect 349342 208046 349398 208102
rect 348970 207922 349026 207978
rect 349094 207922 349150 207978
rect 349218 207922 349274 207978
rect 349342 207922 349398 207978
rect 57250 202294 57306 202350
rect 57374 202294 57430 202350
rect 57498 202294 57554 202350
rect 57622 202294 57678 202350
rect 57250 202170 57306 202226
rect 57374 202170 57430 202226
rect 57498 202170 57554 202226
rect 57622 202170 57678 202226
rect 57250 202046 57306 202102
rect 57374 202046 57430 202102
rect 57498 202046 57554 202102
rect 57622 202046 57678 202102
rect 57250 201922 57306 201978
rect 57374 201922 57430 201978
rect 57498 201922 57554 201978
rect 57622 201922 57678 201978
rect 64518 202294 64574 202350
rect 64642 202294 64698 202350
rect 64518 202170 64574 202226
rect 64642 202170 64698 202226
rect 64518 202046 64574 202102
rect 64642 202046 64698 202102
rect 64518 201922 64574 201978
rect 64642 201922 64698 201978
rect 95238 202294 95294 202350
rect 95362 202294 95418 202350
rect 95238 202170 95294 202226
rect 95362 202170 95418 202226
rect 95238 202046 95294 202102
rect 95362 202046 95418 202102
rect 95238 201922 95294 201978
rect 95362 201922 95418 201978
rect 125958 202294 126014 202350
rect 126082 202294 126138 202350
rect 125958 202170 126014 202226
rect 126082 202170 126138 202226
rect 125958 202046 126014 202102
rect 126082 202046 126138 202102
rect 125958 201922 126014 201978
rect 126082 201922 126138 201978
rect 156678 202294 156734 202350
rect 156802 202294 156858 202350
rect 156678 202170 156734 202226
rect 156802 202170 156858 202226
rect 156678 202046 156734 202102
rect 156802 202046 156858 202102
rect 156678 201922 156734 201978
rect 156802 201922 156858 201978
rect 187398 202294 187454 202350
rect 187522 202294 187578 202350
rect 187398 202170 187454 202226
rect 187522 202170 187578 202226
rect 187398 202046 187454 202102
rect 187522 202046 187578 202102
rect 187398 201922 187454 201978
rect 187522 201922 187578 201978
rect 218118 202294 218174 202350
rect 218242 202294 218298 202350
rect 218118 202170 218174 202226
rect 218242 202170 218298 202226
rect 218118 202046 218174 202102
rect 218242 202046 218298 202102
rect 218118 201922 218174 201978
rect 218242 201922 218298 201978
rect 248838 202294 248894 202350
rect 248962 202294 249018 202350
rect 248838 202170 248894 202226
rect 248962 202170 249018 202226
rect 248838 202046 248894 202102
rect 248962 202046 249018 202102
rect 248838 201922 248894 201978
rect 248962 201922 249018 201978
rect 279558 202294 279614 202350
rect 279682 202294 279738 202350
rect 279558 202170 279614 202226
rect 279682 202170 279738 202226
rect 279558 202046 279614 202102
rect 279682 202046 279738 202102
rect 279558 201922 279614 201978
rect 279682 201922 279738 201978
rect 310278 202294 310334 202350
rect 310402 202294 310458 202350
rect 310278 202170 310334 202226
rect 310402 202170 310458 202226
rect 310278 202046 310334 202102
rect 310402 202046 310458 202102
rect 310278 201922 310334 201978
rect 310402 201922 310458 201978
rect 340998 202294 341054 202350
rect 341122 202294 341178 202350
rect 340998 202170 341054 202226
rect 341122 202170 341178 202226
rect 340998 202046 341054 202102
rect 341122 202046 341178 202102
rect 340998 201922 341054 201978
rect 341122 201922 341178 201978
rect 79878 190294 79934 190350
rect 80002 190294 80058 190350
rect 79878 190170 79934 190226
rect 80002 190170 80058 190226
rect 79878 190046 79934 190102
rect 80002 190046 80058 190102
rect 79878 189922 79934 189978
rect 80002 189922 80058 189978
rect 110598 190294 110654 190350
rect 110722 190294 110778 190350
rect 110598 190170 110654 190226
rect 110722 190170 110778 190226
rect 110598 190046 110654 190102
rect 110722 190046 110778 190102
rect 110598 189922 110654 189978
rect 110722 189922 110778 189978
rect 141318 190294 141374 190350
rect 141442 190294 141498 190350
rect 141318 190170 141374 190226
rect 141442 190170 141498 190226
rect 141318 190046 141374 190102
rect 141442 190046 141498 190102
rect 141318 189922 141374 189978
rect 141442 189922 141498 189978
rect 172038 190294 172094 190350
rect 172162 190294 172218 190350
rect 172038 190170 172094 190226
rect 172162 190170 172218 190226
rect 172038 190046 172094 190102
rect 172162 190046 172218 190102
rect 172038 189922 172094 189978
rect 172162 189922 172218 189978
rect 202758 190294 202814 190350
rect 202882 190294 202938 190350
rect 202758 190170 202814 190226
rect 202882 190170 202938 190226
rect 202758 190046 202814 190102
rect 202882 190046 202938 190102
rect 202758 189922 202814 189978
rect 202882 189922 202938 189978
rect 233478 190294 233534 190350
rect 233602 190294 233658 190350
rect 233478 190170 233534 190226
rect 233602 190170 233658 190226
rect 233478 190046 233534 190102
rect 233602 190046 233658 190102
rect 233478 189922 233534 189978
rect 233602 189922 233658 189978
rect 264198 190294 264254 190350
rect 264322 190294 264378 190350
rect 264198 190170 264254 190226
rect 264322 190170 264378 190226
rect 264198 190046 264254 190102
rect 264322 190046 264378 190102
rect 264198 189922 264254 189978
rect 264322 189922 264378 189978
rect 294918 190294 294974 190350
rect 295042 190294 295098 190350
rect 294918 190170 294974 190226
rect 295042 190170 295098 190226
rect 294918 190046 294974 190102
rect 295042 190046 295098 190102
rect 294918 189922 294974 189978
rect 295042 189922 295098 189978
rect 325638 190294 325694 190350
rect 325762 190294 325818 190350
rect 325638 190170 325694 190226
rect 325762 190170 325818 190226
rect 325638 190046 325694 190102
rect 325762 190046 325818 190102
rect 325638 189922 325694 189978
rect 325762 189922 325818 189978
rect 356358 208294 356414 208350
rect 356482 208294 356538 208350
rect 356358 208170 356414 208226
rect 356482 208170 356538 208226
rect 356358 208046 356414 208102
rect 356482 208046 356538 208102
rect 356358 207922 356414 207978
rect 356482 207922 356538 207978
rect 363250 202294 363306 202350
rect 363374 202294 363430 202350
rect 363498 202294 363554 202350
rect 363622 202294 363678 202350
rect 363250 202170 363306 202226
rect 363374 202170 363430 202226
rect 363498 202170 363554 202226
rect 363622 202170 363678 202226
rect 363250 202046 363306 202102
rect 363374 202046 363430 202102
rect 363498 202046 363554 202102
rect 363622 202046 363678 202102
rect 363250 201922 363306 201978
rect 363374 201922 363430 201978
rect 363498 201922 363554 201978
rect 363622 201922 363678 201978
rect 348970 190294 349026 190350
rect 349094 190294 349150 190350
rect 349218 190294 349274 190350
rect 349342 190294 349398 190350
rect 348970 190170 349026 190226
rect 349094 190170 349150 190226
rect 349218 190170 349274 190226
rect 349342 190170 349398 190226
rect 348970 190046 349026 190102
rect 349094 190046 349150 190102
rect 349218 190046 349274 190102
rect 349342 190046 349398 190102
rect 348970 189922 349026 189978
rect 349094 189922 349150 189978
rect 349218 189922 349274 189978
rect 349342 189922 349398 189978
rect 57250 184294 57306 184350
rect 57374 184294 57430 184350
rect 57498 184294 57554 184350
rect 57622 184294 57678 184350
rect 57250 184170 57306 184226
rect 57374 184170 57430 184226
rect 57498 184170 57554 184226
rect 57622 184170 57678 184226
rect 57250 184046 57306 184102
rect 57374 184046 57430 184102
rect 57498 184046 57554 184102
rect 57622 184046 57678 184102
rect 57250 183922 57306 183978
rect 57374 183922 57430 183978
rect 57498 183922 57554 183978
rect 57622 183922 57678 183978
rect 64518 184294 64574 184350
rect 64642 184294 64698 184350
rect 64518 184170 64574 184226
rect 64642 184170 64698 184226
rect 64518 184046 64574 184102
rect 64642 184046 64698 184102
rect 64518 183922 64574 183978
rect 64642 183922 64698 183978
rect 95238 184294 95294 184350
rect 95362 184294 95418 184350
rect 95238 184170 95294 184226
rect 95362 184170 95418 184226
rect 95238 184046 95294 184102
rect 95362 184046 95418 184102
rect 95238 183922 95294 183978
rect 95362 183922 95418 183978
rect 125958 184294 126014 184350
rect 126082 184294 126138 184350
rect 125958 184170 126014 184226
rect 126082 184170 126138 184226
rect 125958 184046 126014 184102
rect 126082 184046 126138 184102
rect 125958 183922 126014 183978
rect 126082 183922 126138 183978
rect 156678 184294 156734 184350
rect 156802 184294 156858 184350
rect 156678 184170 156734 184226
rect 156802 184170 156858 184226
rect 156678 184046 156734 184102
rect 156802 184046 156858 184102
rect 156678 183922 156734 183978
rect 156802 183922 156858 183978
rect 187398 184294 187454 184350
rect 187522 184294 187578 184350
rect 187398 184170 187454 184226
rect 187522 184170 187578 184226
rect 187398 184046 187454 184102
rect 187522 184046 187578 184102
rect 187398 183922 187454 183978
rect 187522 183922 187578 183978
rect 218118 184294 218174 184350
rect 218242 184294 218298 184350
rect 218118 184170 218174 184226
rect 218242 184170 218298 184226
rect 218118 184046 218174 184102
rect 218242 184046 218298 184102
rect 218118 183922 218174 183978
rect 218242 183922 218298 183978
rect 248838 184294 248894 184350
rect 248962 184294 249018 184350
rect 248838 184170 248894 184226
rect 248962 184170 249018 184226
rect 248838 184046 248894 184102
rect 248962 184046 249018 184102
rect 248838 183922 248894 183978
rect 248962 183922 249018 183978
rect 279558 184294 279614 184350
rect 279682 184294 279738 184350
rect 279558 184170 279614 184226
rect 279682 184170 279738 184226
rect 279558 184046 279614 184102
rect 279682 184046 279738 184102
rect 279558 183922 279614 183978
rect 279682 183922 279738 183978
rect 310278 184294 310334 184350
rect 310402 184294 310458 184350
rect 310278 184170 310334 184226
rect 310402 184170 310458 184226
rect 310278 184046 310334 184102
rect 310402 184046 310458 184102
rect 310278 183922 310334 183978
rect 310402 183922 310458 183978
rect 340998 184294 341054 184350
rect 341122 184294 341178 184350
rect 340998 184170 341054 184226
rect 341122 184170 341178 184226
rect 340998 184046 341054 184102
rect 341122 184046 341178 184102
rect 340998 183922 341054 183978
rect 341122 183922 341178 183978
rect 79878 172294 79934 172350
rect 80002 172294 80058 172350
rect 79878 172170 79934 172226
rect 80002 172170 80058 172226
rect 79878 172046 79934 172102
rect 80002 172046 80058 172102
rect 79878 171922 79934 171978
rect 80002 171922 80058 171978
rect 110598 172294 110654 172350
rect 110722 172294 110778 172350
rect 110598 172170 110654 172226
rect 110722 172170 110778 172226
rect 110598 172046 110654 172102
rect 110722 172046 110778 172102
rect 110598 171922 110654 171978
rect 110722 171922 110778 171978
rect 141318 172294 141374 172350
rect 141442 172294 141498 172350
rect 141318 172170 141374 172226
rect 141442 172170 141498 172226
rect 141318 172046 141374 172102
rect 141442 172046 141498 172102
rect 141318 171922 141374 171978
rect 141442 171922 141498 171978
rect 172038 172294 172094 172350
rect 172162 172294 172218 172350
rect 172038 172170 172094 172226
rect 172162 172170 172218 172226
rect 172038 172046 172094 172102
rect 172162 172046 172218 172102
rect 172038 171922 172094 171978
rect 172162 171922 172218 171978
rect 202758 172294 202814 172350
rect 202882 172294 202938 172350
rect 202758 172170 202814 172226
rect 202882 172170 202938 172226
rect 202758 172046 202814 172102
rect 202882 172046 202938 172102
rect 202758 171922 202814 171978
rect 202882 171922 202938 171978
rect 233478 172294 233534 172350
rect 233602 172294 233658 172350
rect 233478 172170 233534 172226
rect 233602 172170 233658 172226
rect 233478 172046 233534 172102
rect 233602 172046 233658 172102
rect 233478 171922 233534 171978
rect 233602 171922 233658 171978
rect 264198 172294 264254 172350
rect 264322 172294 264378 172350
rect 264198 172170 264254 172226
rect 264322 172170 264378 172226
rect 264198 172046 264254 172102
rect 264322 172046 264378 172102
rect 264198 171922 264254 171978
rect 264322 171922 264378 171978
rect 294918 172294 294974 172350
rect 295042 172294 295098 172350
rect 294918 172170 294974 172226
rect 295042 172170 295098 172226
rect 294918 172046 294974 172102
rect 295042 172046 295098 172102
rect 294918 171922 294974 171978
rect 295042 171922 295098 171978
rect 325638 172294 325694 172350
rect 325762 172294 325818 172350
rect 325638 172170 325694 172226
rect 325762 172170 325818 172226
rect 325638 172046 325694 172102
rect 325762 172046 325818 172102
rect 325638 171922 325694 171978
rect 325762 171922 325818 171978
rect 356358 190294 356414 190350
rect 356482 190294 356538 190350
rect 356358 190170 356414 190226
rect 356482 190170 356538 190226
rect 356358 190046 356414 190102
rect 356482 190046 356538 190102
rect 356358 189922 356414 189978
rect 356482 189922 356538 189978
rect 363250 184294 363306 184350
rect 363374 184294 363430 184350
rect 363498 184294 363554 184350
rect 363622 184294 363678 184350
rect 363250 184170 363306 184226
rect 363374 184170 363430 184226
rect 363498 184170 363554 184226
rect 363622 184170 363678 184226
rect 363250 184046 363306 184102
rect 363374 184046 363430 184102
rect 363498 184046 363554 184102
rect 363622 184046 363678 184102
rect 363250 183922 363306 183978
rect 363374 183922 363430 183978
rect 363498 183922 363554 183978
rect 363622 183922 363678 183978
rect 348970 172294 349026 172350
rect 349094 172294 349150 172350
rect 349218 172294 349274 172350
rect 349342 172294 349398 172350
rect 348970 172170 349026 172226
rect 349094 172170 349150 172226
rect 349218 172170 349274 172226
rect 349342 172170 349398 172226
rect 348970 172046 349026 172102
rect 349094 172046 349150 172102
rect 349218 172046 349274 172102
rect 349342 172046 349398 172102
rect 348970 171922 349026 171978
rect 349094 171922 349150 171978
rect 349218 171922 349274 171978
rect 349342 171922 349398 171978
rect 57250 166294 57306 166350
rect 57374 166294 57430 166350
rect 57498 166294 57554 166350
rect 57622 166294 57678 166350
rect 57250 166170 57306 166226
rect 57374 166170 57430 166226
rect 57498 166170 57554 166226
rect 57622 166170 57678 166226
rect 57250 166046 57306 166102
rect 57374 166046 57430 166102
rect 57498 166046 57554 166102
rect 57622 166046 57678 166102
rect 57250 165922 57306 165978
rect 57374 165922 57430 165978
rect 57498 165922 57554 165978
rect 57622 165922 57678 165978
rect 64518 166294 64574 166350
rect 64642 166294 64698 166350
rect 64518 166170 64574 166226
rect 64642 166170 64698 166226
rect 64518 166046 64574 166102
rect 64642 166046 64698 166102
rect 64518 165922 64574 165978
rect 64642 165922 64698 165978
rect 95238 166294 95294 166350
rect 95362 166294 95418 166350
rect 95238 166170 95294 166226
rect 95362 166170 95418 166226
rect 95238 166046 95294 166102
rect 95362 166046 95418 166102
rect 95238 165922 95294 165978
rect 95362 165922 95418 165978
rect 125958 166294 126014 166350
rect 126082 166294 126138 166350
rect 125958 166170 126014 166226
rect 126082 166170 126138 166226
rect 125958 166046 126014 166102
rect 126082 166046 126138 166102
rect 125958 165922 126014 165978
rect 126082 165922 126138 165978
rect 156678 166294 156734 166350
rect 156802 166294 156858 166350
rect 156678 166170 156734 166226
rect 156802 166170 156858 166226
rect 156678 166046 156734 166102
rect 156802 166046 156858 166102
rect 156678 165922 156734 165978
rect 156802 165922 156858 165978
rect 187398 166294 187454 166350
rect 187522 166294 187578 166350
rect 187398 166170 187454 166226
rect 187522 166170 187578 166226
rect 187398 166046 187454 166102
rect 187522 166046 187578 166102
rect 187398 165922 187454 165978
rect 187522 165922 187578 165978
rect 218118 166294 218174 166350
rect 218242 166294 218298 166350
rect 218118 166170 218174 166226
rect 218242 166170 218298 166226
rect 218118 166046 218174 166102
rect 218242 166046 218298 166102
rect 218118 165922 218174 165978
rect 218242 165922 218298 165978
rect 248838 166294 248894 166350
rect 248962 166294 249018 166350
rect 248838 166170 248894 166226
rect 248962 166170 249018 166226
rect 248838 166046 248894 166102
rect 248962 166046 249018 166102
rect 248838 165922 248894 165978
rect 248962 165922 249018 165978
rect 279558 166294 279614 166350
rect 279682 166294 279738 166350
rect 279558 166170 279614 166226
rect 279682 166170 279738 166226
rect 279558 166046 279614 166102
rect 279682 166046 279738 166102
rect 279558 165922 279614 165978
rect 279682 165922 279738 165978
rect 310278 166294 310334 166350
rect 310402 166294 310458 166350
rect 310278 166170 310334 166226
rect 310402 166170 310458 166226
rect 310278 166046 310334 166102
rect 310402 166046 310458 166102
rect 310278 165922 310334 165978
rect 310402 165922 310458 165978
rect 340998 166294 341054 166350
rect 341122 166294 341178 166350
rect 340998 166170 341054 166226
rect 341122 166170 341178 166226
rect 340998 166046 341054 166102
rect 341122 166046 341178 166102
rect 340998 165922 341054 165978
rect 341122 165922 341178 165978
rect 79878 154294 79934 154350
rect 80002 154294 80058 154350
rect 79878 154170 79934 154226
rect 80002 154170 80058 154226
rect 79878 154046 79934 154102
rect 80002 154046 80058 154102
rect 79878 153922 79934 153978
rect 80002 153922 80058 153978
rect 110598 154294 110654 154350
rect 110722 154294 110778 154350
rect 110598 154170 110654 154226
rect 110722 154170 110778 154226
rect 110598 154046 110654 154102
rect 110722 154046 110778 154102
rect 110598 153922 110654 153978
rect 110722 153922 110778 153978
rect 141318 154294 141374 154350
rect 141442 154294 141498 154350
rect 141318 154170 141374 154226
rect 141442 154170 141498 154226
rect 141318 154046 141374 154102
rect 141442 154046 141498 154102
rect 141318 153922 141374 153978
rect 141442 153922 141498 153978
rect 172038 154294 172094 154350
rect 172162 154294 172218 154350
rect 172038 154170 172094 154226
rect 172162 154170 172218 154226
rect 172038 154046 172094 154102
rect 172162 154046 172218 154102
rect 172038 153922 172094 153978
rect 172162 153922 172218 153978
rect 202758 154294 202814 154350
rect 202882 154294 202938 154350
rect 202758 154170 202814 154226
rect 202882 154170 202938 154226
rect 202758 154046 202814 154102
rect 202882 154046 202938 154102
rect 202758 153922 202814 153978
rect 202882 153922 202938 153978
rect 233478 154294 233534 154350
rect 233602 154294 233658 154350
rect 233478 154170 233534 154226
rect 233602 154170 233658 154226
rect 233478 154046 233534 154102
rect 233602 154046 233658 154102
rect 233478 153922 233534 153978
rect 233602 153922 233658 153978
rect 264198 154294 264254 154350
rect 264322 154294 264378 154350
rect 264198 154170 264254 154226
rect 264322 154170 264378 154226
rect 264198 154046 264254 154102
rect 264322 154046 264378 154102
rect 264198 153922 264254 153978
rect 264322 153922 264378 153978
rect 294918 154294 294974 154350
rect 295042 154294 295098 154350
rect 294918 154170 294974 154226
rect 295042 154170 295098 154226
rect 294918 154046 294974 154102
rect 295042 154046 295098 154102
rect 294918 153922 294974 153978
rect 295042 153922 295098 153978
rect 325638 154294 325694 154350
rect 325762 154294 325818 154350
rect 325638 154170 325694 154226
rect 325762 154170 325818 154226
rect 325638 154046 325694 154102
rect 325762 154046 325818 154102
rect 325638 153922 325694 153978
rect 325762 153922 325818 153978
rect 356358 172294 356414 172350
rect 356482 172294 356538 172350
rect 356358 172170 356414 172226
rect 356482 172170 356538 172226
rect 356358 172046 356414 172102
rect 356482 172046 356538 172102
rect 356358 171922 356414 171978
rect 356482 171922 356538 171978
rect 363250 166294 363306 166350
rect 363374 166294 363430 166350
rect 363498 166294 363554 166350
rect 363622 166294 363678 166350
rect 363250 166170 363306 166226
rect 363374 166170 363430 166226
rect 363498 166170 363554 166226
rect 363622 166170 363678 166226
rect 363250 166046 363306 166102
rect 363374 166046 363430 166102
rect 363498 166046 363554 166102
rect 363622 166046 363678 166102
rect 363250 165922 363306 165978
rect 363374 165922 363430 165978
rect 363498 165922 363554 165978
rect 363622 165922 363678 165978
rect 348970 154294 349026 154350
rect 349094 154294 349150 154350
rect 349218 154294 349274 154350
rect 349342 154294 349398 154350
rect 348970 154170 349026 154226
rect 349094 154170 349150 154226
rect 349218 154170 349274 154226
rect 349342 154170 349398 154226
rect 348970 154046 349026 154102
rect 349094 154046 349150 154102
rect 349218 154046 349274 154102
rect 349342 154046 349398 154102
rect 348970 153922 349026 153978
rect 349094 153922 349150 153978
rect 349218 153922 349274 153978
rect 349342 153922 349398 153978
rect 57250 148294 57306 148350
rect 57374 148294 57430 148350
rect 57498 148294 57554 148350
rect 57622 148294 57678 148350
rect 57250 148170 57306 148226
rect 57374 148170 57430 148226
rect 57498 148170 57554 148226
rect 57622 148170 57678 148226
rect 57250 148046 57306 148102
rect 57374 148046 57430 148102
rect 57498 148046 57554 148102
rect 57622 148046 57678 148102
rect 57250 147922 57306 147978
rect 57374 147922 57430 147978
rect 57498 147922 57554 147978
rect 57622 147922 57678 147978
rect 64518 148294 64574 148350
rect 64642 148294 64698 148350
rect 64518 148170 64574 148226
rect 64642 148170 64698 148226
rect 64518 148046 64574 148102
rect 64642 148046 64698 148102
rect 64518 147922 64574 147978
rect 64642 147922 64698 147978
rect 95238 148294 95294 148350
rect 95362 148294 95418 148350
rect 95238 148170 95294 148226
rect 95362 148170 95418 148226
rect 95238 148046 95294 148102
rect 95362 148046 95418 148102
rect 95238 147922 95294 147978
rect 95362 147922 95418 147978
rect 125958 148294 126014 148350
rect 126082 148294 126138 148350
rect 125958 148170 126014 148226
rect 126082 148170 126138 148226
rect 125958 148046 126014 148102
rect 126082 148046 126138 148102
rect 125958 147922 126014 147978
rect 126082 147922 126138 147978
rect 156678 148294 156734 148350
rect 156802 148294 156858 148350
rect 156678 148170 156734 148226
rect 156802 148170 156858 148226
rect 156678 148046 156734 148102
rect 156802 148046 156858 148102
rect 156678 147922 156734 147978
rect 156802 147922 156858 147978
rect 187398 148294 187454 148350
rect 187522 148294 187578 148350
rect 187398 148170 187454 148226
rect 187522 148170 187578 148226
rect 187398 148046 187454 148102
rect 187522 148046 187578 148102
rect 187398 147922 187454 147978
rect 187522 147922 187578 147978
rect 218118 148294 218174 148350
rect 218242 148294 218298 148350
rect 218118 148170 218174 148226
rect 218242 148170 218298 148226
rect 218118 148046 218174 148102
rect 218242 148046 218298 148102
rect 218118 147922 218174 147978
rect 218242 147922 218298 147978
rect 248838 148294 248894 148350
rect 248962 148294 249018 148350
rect 248838 148170 248894 148226
rect 248962 148170 249018 148226
rect 248838 148046 248894 148102
rect 248962 148046 249018 148102
rect 248838 147922 248894 147978
rect 248962 147922 249018 147978
rect 279558 148294 279614 148350
rect 279682 148294 279738 148350
rect 279558 148170 279614 148226
rect 279682 148170 279738 148226
rect 279558 148046 279614 148102
rect 279682 148046 279738 148102
rect 279558 147922 279614 147978
rect 279682 147922 279738 147978
rect 310278 148294 310334 148350
rect 310402 148294 310458 148350
rect 310278 148170 310334 148226
rect 310402 148170 310458 148226
rect 310278 148046 310334 148102
rect 310402 148046 310458 148102
rect 310278 147922 310334 147978
rect 310402 147922 310458 147978
rect 340998 148294 341054 148350
rect 341122 148294 341178 148350
rect 340998 148170 341054 148226
rect 341122 148170 341178 148226
rect 340998 148046 341054 148102
rect 341122 148046 341178 148102
rect 340998 147922 341054 147978
rect 341122 147922 341178 147978
rect 79878 136294 79934 136350
rect 80002 136294 80058 136350
rect 79878 136170 79934 136226
rect 80002 136170 80058 136226
rect 79878 136046 79934 136102
rect 80002 136046 80058 136102
rect 79878 135922 79934 135978
rect 80002 135922 80058 135978
rect 110598 136294 110654 136350
rect 110722 136294 110778 136350
rect 110598 136170 110654 136226
rect 110722 136170 110778 136226
rect 110598 136046 110654 136102
rect 110722 136046 110778 136102
rect 110598 135922 110654 135978
rect 110722 135922 110778 135978
rect 141318 136294 141374 136350
rect 141442 136294 141498 136350
rect 141318 136170 141374 136226
rect 141442 136170 141498 136226
rect 141318 136046 141374 136102
rect 141442 136046 141498 136102
rect 141318 135922 141374 135978
rect 141442 135922 141498 135978
rect 172038 136294 172094 136350
rect 172162 136294 172218 136350
rect 172038 136170 172094 136226
rect 172162 136170 172218 136226
rect 172038 136046 172094 136102
rect 172162 136046 172218 136102
rect 172038 135922 172094 135978
rect 172162 135922 172218 135978
rect 202758 136294 202814 136350
rect 202882 136294 202938 136350
rect 202758 136170 202814 136226
rect 202882 136170 202938 136226
rect 202758 136046 202814 136102
rect 202882 136046 202938 136102
rect 202758 135922 202814 135978
rect 202882 135922 202938 135978
rect 233478 136294 233534 136350
rect 233602 136294 233658 136350
rect 233478 136170 233534 136226
rect 233602 136170 233658 136226
rect 233478 136046 233534 136102
rect 233602 136046 233658 136102
rect 233478 135922 233534 135978
rect 233602 135922 233658 135978
rect 264198 136294 264254 136350
rect 264322 136294 264378 136350
rect 264198 136170 264254 136226
rect 264322 136170 264378 136226
rect 264198 136046 264254 136102
rect 264322 136046 264378 136102
rect 264198 135922 264254 135978
rect 264322 135922 264378 135978
rect 294918 136294 294974 136350
rect 295042 136294 295098 136350
rect 294918 136170 294974 136226
rect 295042 136170 295098 136226
rect 294918 136046 294974 136102
rect 295042 136046 295098 136102
rect 294918 135922 294974 135978
rect 295042 135922 295098 135978
rect 325638 136294 325694 136350
rect 325762 136294 325818 136350
rect 325638 136170 325694 136226
rect 325762 136170 325818 136226
rect 325638 136046 325694 136102
rect 325762 136046 325818 136102
rect 325638 135922 325694 135978
rect 325762 135922 325818 135978
rect 356358 154294 356414 154350
rect 356482 154294 356538 154350
rect 356358 154170 356414 154226
rect 356482 154170 356538 154226
rect 356358 154046 356414 154102
rect 356482 154046 356538 154102
rect 356358 153922 356414 153978
rect 356482 153922 356538 153978
rect 363250 148294 363306 148350
rect 363374 148294 363430 148350
rect 363498 148294 363554 148350
rect 363622 148294 363678 148350
rect 363250 148170 363306 148226
rect 363374 148170 363430 148226
rect 363498 148170 363554 148226
rect 363622 148170 363678 148226
rect 363250 148046 363306 148102
rect 363374 148046 363430 148102
rect 363498 148046 363554 148102
rect 363622 148046 363678 148102
rect 363250 147922 363306 147978
rect 363374 147922 363430 147978
rect 363498 147922 363554 147978
rect 363622 147922 363678 147978
rect 348970 136294 349026 136350
rect 349094 136294 349150 136350
rect 349218 136294 349274 136350
rect 349342 136294 349398 136350
rect 348970 136170 349026 136226
rect 349094 136170 349150 136226
rect 349218 136170 349274 136226
rect 349342 136170 349398 136226
rect 348970 136046 349026 136102
rect 349094 136046 349150 136102
rect 349218 136046 349274 136102
rect 349342 136046 349398 136102
rect 348970 135922 349026 135978
rect 349094 135922 349150 135978
rect 349218 135922 349274 135978
rect 349342 135922 349398 135978
rect 57250 130294 57306 130350
rect 57374 130294 57430 130350
rect 57498 130294 57554 130350
rect 57622 130294 57678 130350
rect 57250 130170 57306 130226
rect 57374 130170 57430 130226
rect 57498 130170 57554 130226
rect 57622 130170 57678 130226
rect 57250 130046 57306 130102
rect 57374 130046 57430 130102
rect 57498 130046 57554 130102
rect 57622 130046 57678 130102
rect 57250 129922 57306 129978
rect 57374 129922 57430 129978
rect 57498 129922 57554 129978
rect 57622 129922 57678 129978
rect 64518 130294 64574 130350
rect 64642 130294 64698 130350
rect 64518 130170 64574 130226
rect 64642 130170 64698 130226
rect 64518 130046 64574 130102
rect 64642 130046 64698 130102
rect 64518 129922 64574 129978
rect 64642 129922 64698 129978
rect 95238 130294 95294 130350
rect 95362 130294 95418 130350
rect 95238 130170 95294 130226
rect 95362 130170 95418 130226
rect 95238 130046 95294 130102
rect 95362 130046 95418 130102
rect 95238 129922 95294 129978
rect 95362 129922 95418 129978
rect 125958 130294 126014 130350
rect 126082 130294 126138 130350
rect 125958 130170 126014 130226
rect 126082 130170 126138 130226
rect 125958 130046 126014 130102
rect 126082 130046 126138 130102
rect 125958 129922 126014 129978
rect 126082 129922 126138 129978
rect 156678 130294 156734 130350
rect 156802 130294 156858 130350
rect 156678 130170 156734 130226
rect 156802 130170 156858 130226
rect 156678 130046 156734 130102
rect 156802 130046 156858 130102
rect 156678 129922 156734 129978
rect 156802 129922 156858 129978
rect 187398 130294 187454 130350
rect 187522 130294 187578 130350
rect 187398 130170 187454 130226
rect 187522 130170 187578 130226
rect 187398 130046 187454 130102
rect 187522 130046 187578 130102
rect 187398 129922 187454 129978
rect 187522 129922 187578 129978
rect 218118 130294 218174 130350
rect 218242 130294 218298 130350
rect 218118 130170 218174 130226
rect 218242 130170 218298 130226
rect 218118 130046 218174 130102
rect 218242 130046 218298 130102
rect 218118 129922 218174 129978
rect 218242 129922 218298 129978
rect 248838 130294 248894 130350
rect 248962 130294 249018 130350
rect 248838 130170 248894 130226
rect 248962 130170 249018 130226
rect 248838 130046 248894 130102
rect 248962 130046 249018 130102
rect 248838 129922 248894 129978
rect 248962 129922 249018 129978
rect 279558 130294 279614 130350
rect 279682 130294 279738 130350
rect 279558 130170 279614 130226
rect 279682 130170 279738 130226
rect 279558 130046 279614 130102
rect 279682 130046 279738 130102
rect 279558 129922 279614 129978
rect 279682 129922 279738 129978
rect 310278 130294 310334 130350
rect 310402 130294 310458 130350
rect 310278 130170 310334 130226
rect 310402 130170 310458 130226
rect 310278 130046 310334 130102
rect 310402 130046 310458 130102
rect 310278 129922 310334 129978
rect 310402 129922 310458 129978
rect 340998 130294 341054 130350
rect 341122 130294 341178 130350
rect 340998 130170 341054 130226
rect 341122 130170 341178 130226
rect 340998 130046 341054 130102
rect 341122 130046 341178 130102
rect 340998 129922 341054 129978
rect 341122 129922 341178 129978
rect 79878 118294 79934 118350
rect 80002 118294 80058 118350
rect 79878 118170 79934 118226
rect 80002 118170 80058 118226
rect 79878 118046 79934 118102
rect 80002 118046 80058 118102
rect 79878 117922 79934 117978
rect 80002 117922 80058 117978
rect 110598 118294 110654 118350
rect 110722 118294 110778 118350
rect 110598 118170 110654 118226
rect 110722 118170 110778 118226
rect 110598 118046 110654 118102
rect 110722 118046 110778 118102
rect 110598 117922 110654 117978
rect 110722 117922 110778 117978
rect 141318 118294 141374 118350
rect 141442 118294 141498 118350
rect 141318 118170 141374 118226
rect 141442 118170 141498 118226
rect 141318 118046 141374 118102
rect 141442 118046 141498 118102
rect 141318 117922 141374 117978
rect 141442 117922 141498 117978
rect 172038 118294 172094 118350
rect 172162 118294 172218 118350
rect 172038 118170 172094 118226
rect 172162 118170 172218 118226
rect 172038 118046 172094 118102
rect 172162 118046 172218 118102
rect 172038 117922 172094 117978
rect 172162 117922 172218 117978
rect 202758 118294 202814 118350
rect 202882 118294 202938 118350
rect 202758 118170 202814 118226
rect 202882 118170 202938 118226
rect 202758 118046 202814 118102
rect 202882 118046 202938 118102
rect 202758 117922 202814 117978
rect 202882 117922 202938 117978
rect 233478 118294 233534 118350
rect 233602 118294 233658 118350
rect 233478 118170 233534 118226
rect 233602 118170 233658 118226
rect 233478 118046 233534 118102
rect 233602 118046 233658 118102
rect 233478 117922 233534 117978
rect 233602 117922 233658 117978
rect 264198 118294 264254 118350
rect 264322 118294 264378 118350
rect 264198 118170 264254 118226
rect 264322 118170 264378 118226
rect 264198 118046 264254 118102
rect 264322 118046 264378 118102
rect 264198 117922 264254 117978
rect 264322 117922 264378 117978
rect 294918 118294 294974 118350
rect 295042 118294 295098 118350
rect 294918 118170 294974 118226
rect 295042 118170 295098 118226
rect 294918 118046 294974 118102
rect 295042 118046 295098 118102
rect 294918 117922 294974 117978
rect 295042 117922 295098 117978
rect 325638 118294 325694 118350
rect 325762 118294 325818 118350
rect 325638 118170 325694 118226
rect 325762 118170 325818 118226
rect 325638 118046 325694 118102
rect 325762 118046 325818 118102
rect 325638 117922 325694 117978
rect 325762 117922 325818 117978
rect 356358 136294 356414 136350
rect 356482 136294 356538 136350
rect 356358 136170 356414 136226
rect 356482 136170 356538 136226
rect 356358 136046 356414 136102
rect 356482 136046 356538 136102
rect 356358 135922 356414 135978
rect 356482 135922 356538 135978
rect 363250 130294 363306 130350
rect 363374 130294 363430 130350
rect 363498 130294 363554 130350
rect 363622 130294 363678 130350
rect 363250 130170 363306 130226
rect 363374 130170 363430 130226
rect 363498 130170 363554 130226
rect 363622 130170 363678 130226
rect 363250 130046 363306 130102
rect 363374 130046 363430 130102
rect 363498 130046 363554 130102
rect 363622 130046 363678 130102
rect 363250 129922 363306 129978
rect 363374 129922 363430 129978
rect 363498 129922 363554 129978
rect 363622 129922 363678 129978
rect 348970 118294 349026 118350
rect 349094 118294 349150 118350
rect 349218 118294 349274 118350
rect 349342 118294 349398 118350
rect 348970 118170 349026 118226
rect 349094 118170 349150 118226
rect 349218 118170 349274 118226
rect 349342 118170 349398 118226
rect 348970 118046 349026 118102
rect 349094 118046 349150 118102
rect 349218 118046 349274 118102
rect 349342 118046 349398 118102
rect 348970 117922 349026 117978
rect 349094 117922 349150 117978
rect 349218 117922 349274 117978
rect 349342 117922 349398 117978
rect 57250 112294 57306 112350
rect 57374 112294 57430 112350
rect 57498 112294 57554 112350
rect 57622 112294 57678 112350
rect 57250 112170 57306 112226
rect 57374 112170 57430 112226
rect 57498 112170 57554 112226
rect 57622 112170 57678 112226
rect 57250 112046 57306 112102
rect 57374 112046 57430 112102
rect 57498 112046 57554 112102
rect 57622 112046 57678 112102
rect 57250 111922 57306 111978
rect 57374 111922 57430 111978
rect 57498 111922 57554 111978
rect 57622 111922 57678 111978
rect 64518 112294 64574 112350
rect 64642 112294 64698 112350
rect 64518 112170 64574 112226
rect 64642 112170 64698 112226
rect 64518 112046 64574 112102
rect 64642 112046 64698 112102
rect 64518 111922 64574 111978
rect 64642 111922 64698 111978
rect 95238 112294 95294 112350
rect 95362 112294 95418 112350
rect 95238 112170 95294 112226
rect 95362 112170 95418 112226
rect 95238 112046 95294 112102
rect 95362 112046 95418 112102
rect 95238 111922 95294 111978
rect 95362 111922 95418 111978
rect 125958 112294 126014 112350
rect 126082 112294 126138 112350
rect 125958 112170 126014 112226
rect 126082 112170 126138 112226
rect 125958 112046 126014 112102
rect 126082 112046 126138 112102
rect 125958 111922 126014 111978
rect 126082 111922 126138 111978
rect 156678 112294 156734 112350
rect 156802 112294 156858 112350
rect 156678 112170 156734 112226
rect 156802 112170 156858 112226
rect 156678 112046 156734 112102
rect 156802 112046 156858 112102
rect 156678 111922 156734 111978
rect 156802 111922 156858 111978
rect 187398 112294 187454 112350
rect 187522 112294 187578 112350
rect 187398 112170 187454 112226
rect 187522 112170 187578 112226
rect 187398 112046 187454 112102
rect 187522 112046 187578 112102
rect 187398 111922 187454 111978
rect 187522 111922 187578 111978
rect 218118 112294 218174 112350
rect 218242 112294 218298 112350
rect 218118 112170 218174 112226
rect 218242 112170 218298 112226
rect 218118 112046 218174 112102
rect 218242 112046 218298 112102
rect 218118 111922 218174 111978
rect 218242 111922 218298 111978
rect 248838 112294 248894 112350
rect 248962 112294 249018 112350
rect 248838 112170 248894 112226
rect 248962 112170 249018 112226
rect 248838 112046 248894 112102
rect 248962 112046 249018 112102
rect 248838 111922 248894 111978
rect 248962 111922 249018 111978
rect 279558 112294 279614 112350
rect 279682 112294 279738 112350
rect 279558 112170 279614 112226
rect 279682 112170 279738 112226
rect 279558 112046 279614 112102
rect 279682 112046 279738 112102
rect 279558 111922 279614 111978
rect 279682 111922 279738 111978
rect 310278 112294 310334 112350
rect 310402 112294 310458 112350
rect 310278 112170 310334 112226
rect 310402 112170 310458 112226
rect 310278 112046 310334 112102
rect 310402 112046 310458 112102
rect 310278 111922 310334 111978
rect 310402 111922 310458 111978
rect 340998 112294 341054 112350
rect 341122 112294 341178 112350
rect 340998 112170 341054 112226
rect 341122 112170 341178 112226
rect 340998 112046 341054 112102
rect 341122 112046 341178 112102
rect 340998 111922 341054 111978
rect 341122 111922 341178 111978
rect 79878 100294 79934 100350
rect 80002 100294 80058 100350
rect 79878 100170 79934 100226
rect 80002 100170 80058 100226
rect 79878 100046 79934 100102
rect 80002 100046 80058 100102
rect 79878 99922 79934 99978
rect 80002 99922 80058 99978
rect 110598 100294 110654 100350
rect 110722 100294 110778 100350
rect 110598 100170 110654 100226
rect 110722 100170 110778 100226
rect 110598 100046 110654 100102
rect 110722 100046 110778 100102
rect 110598 99922 110654 99978
rect 110722 99922 110778 99978
rect 141318 100294 141374 100350
rect 141442 100294 141498 100350
rect 141318 100170 141374 100226
rect 141442 100170 141498 100226
rect 141318 100046 141374 100102
rect 141442 100046 141498 100102
rect 141318 99922 141374 99978
rect 141442 99922 141498 99978
rect 172038 100294 172094 100350
rect 172162 100294 172218 100350
rect 172038 100170 172094 100226
rect 172162 100170 172218 100226
rect 172038 100046 172094 100102
rect 172162 100046 172218 100102
rect 172038 99922 172094 99978
rect 172162 99922 172218 99978
rect 202758 100294 202814 100350
rect 202882 100294 202938 100350
rect 202758 100170 202814 100226
rect 202882 100170 202938 100226
rect 202758 100046 202814 100102
rect 202882 100046 202938 100102
rect 202758 99922 202814 99978
rect 202882 99922 202938 99978
rect 233478 100294 233534 100350
rect 233602 100294 233658 100350
rect 233478 100170 233534 100226
rect 233602 100170 233658 100226
rect 233478 100046 233534 100102
rect 233602 100046 233658 100102
rect 233478 99922 233534 99978
rect 233602 99922 233658 99978
rect 264198 100294 264254 100350
rect 264322 100294 264378 100350
rect 264198 100170 264254 100226
rect 264322 100170 264378 100226
rect 264198 100046 264254 100102
rect 264322 100046 264378 100102
rect 264198 99922 264254 99978
rect 264322 99922 264378 99978
rect 294918 100294 294974 100350
rect 295042 100294 295098 100350
rect 294918 100170 294974 100226
rect 295042 100170 295098 100226
rect 294918 100046 294974 100102
rect 295042 100046 295098 100102
rect 294918 99922 294974 99978
rect 295042 99922 295098 99978
rect 325638 100294 325694 100350
rect 325762 100294 325818 100350
rect 325638 100170 325694 100226
rect 325762 100170 325818 100226
rect 325638 100046 325694 100102
rect 325762 100046 325818 100102
rect 325638 99922 325694 99978
rect 325762 99922 325818 99978
rect 356358 118294 356414 118350
rect 356482 118294 356538 118350
rect 356358 118170 356414 118226
rect 356482 118170 356538 118226
rect 356358 118046 356414 118102
rect 356482 118046 356538 118102
rect 356358 117922 356414 117978
rect 356482 117922 356538 117978
rect 363250 112294 363306 112350
rect 363374 112294 363430 112350
rect 363498 112294 363554 112350
rect 363622 112294 363678 112350
rect 363250 112170 363306 112226
rect 363374 112170 363430 112226
rect 363498 112170 363554 112226
rect 363622 112170 363678 112226
rect 363250 112046 363306 112102
rect 363374 112046 363430 112102
rect 363498 112046 363554 112102
rect 363622 112046 363678 112102
rect 363250 111922 363306 111978
rect 363374 111922 363430 111978
rect 363498 111922 363554 111978
rect 363622 111922 363678 111978
rect 348970 100294 349026 100350
rect 349094 100294 349150 100350
rect 349218 100294 349274 100350
rect 349342 100294 349398 100350
rect 348970 100170 349026 100226
rect 349094 100170 349150 100226
rect 349218 100170 349274 100226
rect 349342 100170 349398 100226
rect 348970 100046 349026 100102
rect 349094 100046 349150 100102
rect 349218 100046 349274 100102
rect 349342 100046 349398 100102
rect 348970 99922 349026 99978
rect 349094 99922 349150 99978
rect 349218 99922 349274 99978
rect 349342 99922 349398 99978
rect 57250 94294 57306 94350
rect 57374 94294 57430 94350
rect 57498 94294 57554 94350
rect 57622 94294 57678 94350
rect 57250 94170 57306 94226
rect 57374 94170 57430 94226
rect 57498 94170 57554 94226
rect 57622 94170 57678 94226
rect 57250 94046 57306 94102
rect 57374 94046 57430 94102
rect 57498 94046 57554 94102
rect 57622 94046 57678 94102
rect 57250 93922 57306 93978
rect 57374 93922 57430 93978
rect 57498 93922 57554 93978
rect 57622 93922 57678 93978
rect 64518 94294 64574 94350
rect 64642 94294 64698 94350
rect 64518 94170 64574 94226
rect 64642 94170 64698 94226
rect 64518 94046 64574 94102
rect 64642 94046 64698 94102
rect 64518 93922 64574 93978
rect 64642 93922 64698 93978
rect 95238 94294 95294 94350
rect 95362 94294 95418 94350
rect 95238 94170 95294 94226
rect 95362 94170 95418 94226
rect 95238 94046 95294 94102
rect 95362 94046 95418 94102
rect 95238 93922 95294 93978
rect 95362 93922 95418 93978
rect 125958 94294 126014 94350
rect 126082 94294 126138 94350
rect 125958 94170 126014 94226
rect 126082 94170 126138 94226
rect 125958 94046 126014 94102
rect 126082 94046 126138 94102
rect 125958 93922 126014 93978
rect 126082 93922 126138 93978
rect 156678 94294 156734 94350
rect 156802 94294 156858 94350
rect 156678 94170 156734 94226
rect 156802 94170 156858 94226
rect 156678 94046 156734 94102
rect 156802 94046 156858 94102
rect 156678 93922 156734 93978
rect 156802 93922 156858 93978
rect 187398 94294 187454 94350
rect 187522 94294 187578 94350
rect 187398 94170 187454 94226
rect 187522 94170 187578 94226
rect 187398 94046 187454 94102
rect 187522 94046 187578 94102
rect 187398 93922 187454 93978
rect 187522 93922 187578 93978
rect 218118 94294 218174 94350
rect 218242 94294 218298 94350
rect 218118 94170 218174 94226
rect 218242 94170 218298 94226
rect 218118 94046 218174 94102
rect 218242 94046 218298 94102
rect 218118 93922 218174 93978
rect 218242 93922 218298 93978
rect 248838 94294 248894 94350
rect 248962 94294 249018 94350
rect 248838 94170 248894 94226
rect 248962 94170 249018 94226
rect 248838 94046 248894 94102
rect 248962 94046 249018 94102
rect 248838 93922 248894 93978
rect 248962 93922 249018 93978
rect 279558 94294 279614 94350
rect 279682 94294 279738 94350
rect 279558 94170 279614 94226
rect 279682 94170 279738 94226
rect 279558 94046 279614 94102
rect 279682 94046 279738 94102
rect 279558 93922 279614 93978
rect 279682 93922 279738 93978
rect 310278 94294 310334 94350
rect 310402 94294 310458 94350
rect 310278 94170 310334 94226
rect 310402 94170 310458 94226
rect 310278 94046 310334 94102
rect 310402 94046 310458 94102
rect 310278 93922 310334 93978
rect 310402 93922 310458 93978
rect 340998 94294 341054 94350
rect 341122 94294 341178 94350
rect 340998 94170 341054 94226
rect 341122 94170 341178 94226
rect 340998 94046 341054 94102
rect 341122 94046 341178 94102
rect 340998 93922 341054 93978
rect 341122 93922 341178 93978
rect 79878 82294 79934 82350
rect 80002 82294 80058 82350
rect 79878 82170 79934 82226
rect 80002 82170 80058 82226
rect 79878 82046 79934 82102
rect 80002 82046 80058 82102
rect 79878 81922 79934 81978
rect 80002 81922 80058 81978
rect 110598 82294 110654 82350
rect 110722 82294 110778 82350
rect 110598 82170 110654 82226
rect 110722 82170 110778 82226
rect 110598 82046 110654 82102
rect 110722 82046 110778 82102
rect 110598 81922 110654 81978
rect 110722 81922 110778 81978
rect 141318 82294 141374 82350
rect 141442 82294 141498 82350
rect 141318 82170 141374 82226
rect 141442 82170 141498 82226
rect 141318 82046 141374 82102
rect 141442 82046 141498 82102
rect 141318 81922 141374 81978
rect 141442 81922 141498 81978
rect 172038 82294 172094 82350
rect 172162 82294 172218 82350
rect 172038 82170 172094 82226
rect 172162 82170 172218 82226
rect 172038 82046 172094 82102
rect 172162 82046 172218 82102
rect 172038 81922 172094 81978
rect 172162 81922 172218 81978
rect 202758 82294 202814 82350
rect 202882 82294 202938 82350
rect 202758 82170 202814 82226
rect 202882 82170 202938 82226
rect 202758 82046 202814 82102
rect 202882 82046 202938 82102
rect 202758 81922 202814 81978
rect 202882 81922 202938 81978
rect 233478 82294 233534 82350
rect 233602 82294 233658 82350
rect 233478 82170 233534 82226
rect 233602 82170 233658 82226
rect 233478 82046 233534 82102
rect 233602 82046 233658 82102
rect 233478 81922 233534 81978
rect 233602 81922 233658 81978
rect 264198 82294 264254 82350
rect 264322 82294 264378 82350
rect 264198 82170 264254 82226
rect 264322 82170 264378 82226
rect 264198 82046 264254 82102
rect 264322 82046 264378 82102
rect 264198 81922 264254 81978
rect 264322 81922 264378 81978
rect 294918 82294 294974 82350
rect 295042 82294 295098 82350
rect 294918 82170 294974 82226
rect 295042 82170 295098 82226
rect 294918 82046 294974 82102
rect 295042 82046 295098 82102
rect 294918 81922 294974 81978
rect 295042 81922 295098 81978
rect 325638 82294 325694 82350
rect 325762 82294 325818 82350
rect 325638 82170 325694 82226
rect 325762 82170 325818 82226
rect 325638 82046 325694 82102
rect 325762 82046 325818 82102
rect 325638 81922 325694 81978
rect 325762 81922 325818 81978
rect 356358 100294 356414 100350
rect 356482 100294 356538 100350
rect 356358 100170 356414 100226
rect 356482 100170 356538 100226
rect 356358 100046 356414 100102
rect 356482 100046 356538 100102
rect 356358 99922 356414 99978
rect 356482 99922 356538 99978
rect 363250 94294 363306 94350
rect 363374 94294 363430 94350
rect 363498 94294 363554 94350
rect 363622 94294 363678 94350
rect 363250 94170 363306 94226
rect 363374 94170 363430 94226
rect 363498 94170 363554 94226
rect 363622 94170 363678 94226
rect 363250 94046 363306 94102
rect 363374 94046 363430 94102
rect 363498 94046 363554 94102
rect 363622 94046 363678 94102
rect 363250 93922 363306 93978
rect 363374 93922 363430 93978
rect 363498 93922 363554 93978
rect 363622 93922 363678 93978
rect 348970 82294 349026 82350
rect 349094 82294 349150 82350
rect 349218 82294 349274 82350
rect 349342 82294 349398 82350
rect 348970 82170 349026 82226
rect 349094 82170 349150 82226
rect 349218 82170 349274 82226
rect 349342 82170 349398 82226
rect 348970 82046 349026 82102
rect 349094 82046 349150 82102
rect 349218 82046 349274 82102
rect 349342 82046 349398 82102
rect 348970 81922 349026 81978
rect 349094 81922 349150 81978
rect 349218 81922 349274 81978
rect 349342 81922 349398 81978
rect 57250 76294 57306 76350
rect 57374 76294 57430 76350
rect 57498 76294 57554 76350
rect 57622 76294 57678 76350
rect 57250 76170 57306 76226
rect 57374 76170 57430 76226
rect 57498 76170 57554 76226
rect 57622 76170 57678 76226
rect 57250 76046 57306 76102
rect 57374 76046 57430 76102
rect 57498 76046 57554 76102
rect 57622 76046 57678 76102
rect 57250 75922 57306 75978
rect 57374 75922 57430 75978
rect 57498 75922 57554 75978
rect 57622 75922 57678 75978
rect 64518 76294 64574 76350
rect 64642 76294 64698 76350
rect 64518 76170 64574 76226
rect 64642 76170 64698 76226
rect 64518 76046 64574 76102
rect 64642 76046 64698 76102
rect 64518 75922 64574 75978
rect 64642 75922 64698 75978
rect 95238 76294 95294 76350
rect 95362 76294 95418 76350
rect 95238 76170 95294 76226
rect 95362 76170 95418 76226
rect 95238 76046 95294 76102
rect 95362 76046 95418 76102
rect 95238 75922 95294 75978
rect 95362 75922 95418 75978
rect 125958 76294 126014 76350
rect 126082 76294 126138 76350
rect 125958 76170 126014 76226
rect 126082 76170 126138 76226
rect 125958 76046 126014 76102
rect 126082 76046 126138 76102
rect 125958 75922 126014 75978
rect 126082 75922 126138 75978
rect 156678 76294 156734 76350
rect 156802 76294 156858 76350
rect 156678 76170 156734 76226
rect 156802 76170 156858 76226
rect 156678 76046 156734 76102
rect 156802 76046 156858 76102
rect 156678 75922 156734 75978
rect 156802 75922 156858 75978
rect 187398 76294 187454 76350
rect 187522 76294 187578 76350
rect 187398 76170 187454 76226
rect 187522 76170 187578 76226
rect 187398 76046 187454 76102
rect 187522 76046 187578 76102
rect 187398 75922 187454 75978
rect 187522 75922 187578 75978
rect 218118 76294 218174 76350
rect 218242 76294 218298 76350
rect 218118 76170 218174 76226
rect 218242 76170 218298 76226
rect 218118 76046 218174 76102
rect 218242 76046 218298 76102
rect 218118 75922 218174 75978
rect 218242 75922 218298 75978
rect 248838 76294 248894 76350
rect 248962 76294 249018 76350
rect 248838 76170 248894 76226
rect 248962 76170 249018 76226
rect 248838 76046 248894 76102
rect 248962 76046 249018 76102
rect 248838 75922 248894 75978
rect 248962 75922 249018 75978
rect 279558 76294 279614 76350
rect 279682 76294 279738 76350
rect 279558 76170 279614 76226
rect 279682 76170 279738 76226
rect 279558 76046 279614 76102
rect 279682 76046 279738 76102
rect 279558 75922 279614 75978
rect 279682 75922 279738 75978
rect 310278 76294 310334 76350
rect 310402 76294 310458 76350
rect 310278 76170 310334 76226
rect 310402 76170 310458 76226
rect 310278 76046 310334 76102
rect 310402 76046 310458 76102
rect 310278 75922 310334 75978
rect 310402 75922 310458 75978
rect 340998 76294 341054 76350
rect 341122 76294 341178 76350
rect 340998 76170 341054 76226
rect 341122 76170 341178 76226
rect 340998 76046 341054 76102
rect 341122 76046 341178 76102
rect 340998 75922 341054 75978
rect 341122 75922 341178 75978
rect 79878 64294 79934 64350
rect 80002 64294 80058 64350
rect 79878 64170 79934 64226
rect 80002 64170 80058 64226
rect 79878 64046 79934 64102
rect 80002 64046 80058 64102
rect 79878 63922 79934 63978
rect 80002 63922 80058 63978
rect 110598 64294 110654 64350
rect 110722 64294 110778 64350
rect 110598 64170 110654 64226
rect 110722 64170 110778 64226
rect 110598 64046 110654 64102
rect 110722 64046 110778 64102
rect 110598 63922 110654 63978
rect 110722 63922 110778 63978
rect 141318 64294 141374 64350
rect 141442 64294 141498 64350
rect 141318 64170 141374 64226
rect 141442 64170 141498 64226
rect 141318 64046 141374 64102
rect 141442 64046 141498 64102
rect 141318 63922 141374 63978
rect 141442 63922 141498 63978
rect 172038 64294 172094 64350
rect 172162 64294 172218 64350
rect 172038 64170 172094 64226
rect 172162 64170 172218 64226
rect 172038 64046 172094 64102
rect 172162 64046 172218 64102
rect 172038 63922 172094 63978
rect 172162 63922 172218 63978
rect 202758 64294 202814 64350
rect 202882 64294 202938 64350
rect 202758 64170 202814 64226
rect 202882 64170 202938 64226
rect 202758 64046 202814 64102
rect 202882 64046 202938 64102
rect 202758 63922 202814 63978
rect 202882 63922 202938 63978
rect 233478 64294 233534 64350
rect 233602 64294 233658 64350
rect 233478 64170 233534 64226
rect 233602 64170 233658 64226
rect 233478 64046 233534 64102
rect 233602 64046 233658 64102
rect 233478 63922 233534 63978
rect 233602 63922 233658 63978
rect 264198 64294 264254 64350
rect 264322 64294 264378 64350
rect 264198 64170 264254 64226
rect 264322 64170 264378 64226
rect 264198 64046 264254 64102
rect 264322 64046 264378 64102
rect 264198 63922 264254 63978
rect 264322 63922 264378 63978
rect 294918 64294 294974 64350
rect 295042 64294 295098 64350
rect 294918 64170 294974 64226
rect 295042 64170 295098 64226
rect 294918 64046 294974 64102
rect 295042 64046 295098 64102
rect 294918 63922 294974 63978
rect 295042 63922 295098 63978
rect 325638 64294 325694 64350
rect 325762 64294 325818 64350
rect 325638 64170 325694 64226
rect 325762 64170 325818 64226
rect 325638 64046 325694 64102
rect 325762 64046 325818 64102
rect 325638 63922 325694 63978
rect 325762 63922 325818 63978
rect 356358 82294 356414 82350
rect 356482 82294 356538 82350
rect 356358 82170 356414 82226
rect 356482 82170 356538 82226
rect 356358 82046 356414 82102
rect 356482 82046 356538 82102
rect 356358 81922 356414 81978
rect 356482 81922 356538 81978
rect 363250 76294 363306 76350
rect 363374 76294 363430 76350
rect 363498 76294 363554 76350
rect 363622 76294 363678 76350
rect 363250 76170 363306 76226
rect 363374 76170 363430 76226
rect 363498 76170 363554 76226
rect 363622 76170 363678 76226
rect 363250 76046 363306 76102
rect 363374 76046 363430 76102
rect 363498 76046 363554 76102
rect 363622 76046 363678 76102
rect 363250 75922 363306 75978
rect 363374 75922 363430 75978
rect 363498 75922 363554 75978
rect 363622 75922 363678 75978
rect 348970 64294 349026 64350
rect 349094 64294 349150 64350
rect 349218 64294 349274 64350
rect 349342 64294 349398 64350
rect 348970 64170 349026 64226
rect 349094 64170 349150 64226
rect 349218 64170 349274 64226
rect 349342 64170 349398 64226
rect 348970 64046 349026 64102
rect 349094 64046 349150 64102
rect 349218 64046 349274 64102
rect 349342 64046 349398 64102
rect 348970 63922 349026 63978
rect 349094 63922 349150 63978
rect 349218 63922 349274 63978
rect 349342 63922 349398 63978
rect 57250 58294 57306 58350
rect 57374 58294 57430 58350
rect 57498 58294 57554 58350
rect 57622 58294 57678 58350
rect 57250 58170 57306 58226
rect 57374 58170 57430 58226
rect 57498 58170 57554 58226
rect 57622 58170 57678 58226
rect 57250 58046 57306 58102
rect 57374 58046 57430 58102
rect 57498 58046 57554 58102
rect 57622 58046 57678 58102
rect 57250 57922 57306 57978
rect 57374 57922 57430 57978
rect 57498 57922 57554 57978
rect 57622 57922 57678 57978
rect 57250 40294 57306 40350
rect 57374 40294 57430 40350
rect 57498 40294 57554 40350
rect 57622 40294 57678 40350
rect 57250 40170 57306 40226
rect 57374 40170 57430 40226
rect 57498 40170 57554 40226
rect 57622 40170 57678 40226
rect 57250 40046 57306 40102
rect 57374 40046 57430 40102
rect 57498 40046 57554 40102
rect 57622 40046 57678 40102
rect 57250 39922 57306 39978
rect 57374 39922 57430 39978
rect 57498 39922 57554 39978
rect 57622 39922 57678 39978
rect 57250 22294 57306 22350
rect 57374 22294 57430 22350
rect 57498 22294 57554 22350
rect 57622 22294 57678 22350
rect 57250 22170 57306 22226
rect 57374 22170 57430 22226
rect 57498 22170 57554 22226
rect 57622 22170 57678 22226
rect 57250 22046 57306 22102
rect 57374 22046 57430 22102
rect 57498 22046 57554 22102
rect 57622 22046 57678 22102
rect 57250 21922 57306 21978
rect 57374 21922 57430 21978
rect 57498 21922 57554 21978
rect 57622 21922 57678 21978
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 60970 46294 61026 46350
rect 61094 46294 61150 46350
rect 61218 46294 61274 46350
rect 61342 46294 61398 46350
rect 60970 46170 61026 46226
rect 61094 46170 61150 46226
rect 61218 46170 61274 46226
rect 61342 46170 61398 46226
rect 60970 46046 61026 46102
rect 61094 46046 61150 46102
rect 61218 46046 61274 46102
rect 61342 46046 61398 46102
rect 60970 45922 61026 45978
rect 61094 45922 61150 45978
rect 61218 45922 61274 45978
rect 61342 45922 61398 45978
rect 60970 28294 61026 28350
rect 61094 28294 61150 28350
rect 61218 28294 61274 28350
rect 61342 28294 61398 28350
rect 60970 28170 61026 28226
rect 61094 28170 61150 28226
rect 61218 28170 61274 28226
rect 61342 28170 61398 28226
rect 60970 28046 61026 28102
rect 61094 28046 61150 28102
rect 61218 28046 61274 28102
rect 61342 28046 61398 28102
rect 60970 27922 61026 27978
rect 61094 27922 61150 27978
rect 61218 27922 61274 27978
rect 61342 27922 61398 27978
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 58294 75306 58350
rect 75374 58294 75430 58350
rect 75498 58294 75554 58350
rect 75622 58294 75678 58350
rect 75250 58170 75306 58226
rect 75374 58170 75430 58226
rect 75498 58170 75554 58226
rect 75622 58170 75678 58226
rect 75250 58046 75306 58102
rect 75374 58046 75430 58102
rect 75498 58046 75554 58102
rect 75622 58046 75678 58102
rect 75250 57922 75306 57978
rect 75374 57922 75430 57978
rect 75498 57922 75554 57978
rect 75622 57922 75678 57978
rect 75250 40294 75306 40350
rect 75374 40294 75430 40350
rect 75498 40294 75554 40350
rect 75622 40294 75678 40350
rect 75250 40170 75306 40226
rect 75374 40170 75430 40226
rect 75498 40170 75554 40226
rect 75622 40170 75678 40226
rect 75250 40046 75306 40102
rect 75374 40046 75430 40102
rect 75498 40046 75554 40102
rect 75622 40046 75678 40102
rect 75250 39922 75306 39978
rect 75374 39922 75430 39978
rect 75498 39922 75554 39978
rect 75622 39922 75678 39978
rect 75250 22294 75306 22350
rect 75374 22294 75430 22350
rect 75498 22294 75554 22350
rect 75622 22294 75678 22350
rect 75250 22170 75306 22226
rect 75374 22170 75430 22226
rect 75498 22170 75554 22226
rect 75622 22170 75678 22226
rect 75250 22046 75306 22102
rect 75374 22046 75430 22102
rect 75498 22046 75554 22102
rect 75622 22046 75678 22102
rect 75250 21922 75306 21978
rect 75374 21922 75430 21978
rect 75498 21922 75554 21978
rect 75622 21922 75678 21978
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 46294 79026 46350
rect 79094 46294 79150 46350
rect 79218 46294 79274 46350
rect 79342 46294 79398 46350
rect 78970 46170 79026 46226
rect 79094 46170 79150 46226
rect 79218 46170 79274 46226
rect 79342 46170 79398 46226
rect 78970 46046 79026 46102
rect 79094 46046 79150 46102
rect 79218 46046 79274 46102
rect 79342 46046 79398 46102
rect 78970 45922 79026 45978
rect 79094 45922 79150 45978
rect 79218 45922 79274 45978
rect 79342 45922 79398 45978
rect 78970 28294 79026 28350
rect 79094 28294 79150 28350
rect 79218 28294 79274 28350
rect 79342 28294 79398 28350
rect 78970 28170 79026 28226
rect 79094 28170 79150 28226
rect 79218 28170 79274 28226
rect 79342 28170 79398 28226
rect 78970 28046 79026 28102
rect 79094 28046 79150 28102
rect 79218 28046 79274 28102
rect 79342 28046 79398 28102
rect 78970 27922 79026 27978
rect 79094 27922 79150 27978
rect 79218 27922 79274 27978
rect 79342 27922 79398 27978
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 58294 93306 58350
rect 93374 58294 93430 58350
rect 93498 58294 93554 58350
rect 93622 58294 93678 58350
rect 93250 58170 93306 58226
rect 93374 58170 93430 58226
rect 93498 58170 93554 58226
rect 93622 58170 93678 58226
rect 93250 58046 93306 58102
rect 93374 58046 93430 58102
rect 93498 58046 93554 58102
rect 93622 58046 93678 58102
rect 93250 57922 93306 57978
rect 93374 57922 93430 57978
rect 93498 57922 93554 57978
rect 93622 57922 93678 57978
rect 93250 40294 93306 40350
rect 93374 40294 93430 40350
rect 93498 40294 93554 40350
rect 93622 40294 93678 40350
rect 93250 40170 93306 40226
rect 93374 40170 93430 40226
rect 93498 40170 93554 40226
rect 93622 40170 93678 40226
rect 93250 40046 93306 40102
rect 93374 40046 93430 40102
rect 93498 40046 93554 40102
rect 93622 40046 93678 40102
rect 93250 39922 93306 39978
rect 93374 39922 93430 39978
rect 93498 39922 93554 39978
rect 93622 39922 93678 39978
rect 93250 22294 93306 22350
rect 93374 22294 93430 22350
rect 93498 22294 93554 22350
rect 93622 22294 93678 22350
rect 93250 22170 93306 22226
rect 93374 22170 93430 22226
rect 93498 22170 93554 22226
rect 93622 22170 93678 22226
rect 93250 22046 93306 22102
rect 93374 22046 93430 22102
rect 93498 22046 93554 22102
rect 93622 22046 93678 22102
rect 93250 21922 93306 21978
rect 93374 21922 93430 21978
rect 93498 21922 93554 21978
rect 93622 21922 93678 21978
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 96970 46294 97026 46350
rect 97094 46294 97150 46350
rect 97218 46294 97274 46350
rect 97342 46294 97398 46350
rect 96970 46170 97026 46226
rect 97094 46170 97150 46226
rect 97218 46170 97274 46226
rect 97342 46170 97398 46226
rect 96970 46046 97026 46102
rect 97094 46046 97150 46102
rect 97218 46046 97274 46102
rect 97342 46046 97398 46102
rect 96970 45922 97026 45978
rect 97094 45922 97150 45978
rect 97218 45922 97274 45978
rect 97342 45922 97398 45978
rect 96970 28294 97026 28350
rect 97094 28294 97150 28350
rect 97218 28294 97274 28350
rect 97342 28294 97398 28350
rect 96970 28170 97026 28226
rect 97094 28170 97150 28226
rect 97218 28170 97274 28226
rect 97342 28170 97398 28226
rect 96970 28046 97026 28102
rect 97094 28046 97150 28102
rect 97218 28046 97274 28102
rect 97342 28046 97398 28102
rect 96970 27922 97026 27978
rect 97094 27922 97150 27978
rect 97218 27922 97274 27978
rect 97342 27922 97398 27978
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 111250 58294 111306 58350
rect 111374 58294 111430 58350
rect 111498 58294 111554 58350
rect 111622 58294 111678 58350
rect 111250 58170 111306 58226
rect 111374 58170 111430 58226
rect 111498 58170 111554 58226
rect 111622 58170 111678 58226
rect 111250 58046 111306 58102
rect 111374 58046 111430 58102
rect 111498 58046 111554 58102
rect 111622 58046 111678 58102
rect 111250 57922 111306 57978
rect 111374 57922 111430 57978
rect 111498 57922 111554 57978
rect 111622 57922 111678 57978
rect 111250 40294 111306 40350
rect 111374 40294 111430 40350
rect 111498 40294 111554 40350
rect 111622 40294 111678 40350
rect 111250 40170 111306 40226
rect 111374 40170 111430 40226
rect 111498 40170 111554 40226
rect 111622 40170 111678 40226
rect 111250 40046 111306 40102
rect 111374 40046 111430 40102
rect 111498 40046 111554 40102
rect 111622 40046 111678 40102
rect 111250 39922 111306 39978
rect 111374 39922 111430 39978
rect 111498 39922 111554 39978
rect 111622 39922 111678 39978
rect 111250 22294 111306 22350
rect 111374 22294 111430 22350
rect 111498 22294 111554 22350
rect 111622 22294 111678 22350
rect 111250 22170 111306 22226
rect 111374 22170 111430 22226
rect 111498 22170 111554 22226
rect 111622 22170 111678 22226
rect 111250 22046 111306 22102
rect 111374 22046 111430 22102
rect 111498 22046 111554 22102
rect 111622 22046 111678 22102
rect 111250 21922 111306 21978
rect 111374 21922 111430 21978
rect 111498 21922 111554 21978
rect 111622 21922 111678 21978
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 46294 115026 46350
rect 115094 46294 115150 46350
rect 115218 46294 115274 46350
rect 115342 46294 115398 46350
rect 114970 46170 115026 46226
rect 115094 46170 115150 46226
rect 115218 46170 115274 46226
rect 115342 46170 115398 46226
rect 114970 46046 115026 46102
rect 115094 46046 115150 46102
rect 115218 46046 115274 46102
rect 115342 46046 115398 46102
rect 114970 45922 115026 45978
rect 115094 45922 115150 45978
rect 115218 45922 115274 45978
rect 115342 45922 115398 45978
rect 114970 28294 115026 28350
rect 115094 28294 115150 28350
rect 115218 28294 115274 28350
rect 115342 28294 115398 28350
rect 114970 28170 115026 28226
rect 115094 28170 115150 28226
rect 115218 28170 115274 28226
rect 115342 28170 115398 28226
rect 114970 28046 115026 28102
rect 115094 28046 115150 28102
rect 115218 28046 115274 28102
rect 115342 28046 115398 28102
rect 114970 27922 115026 27978
rect 115094 27922 115150 27978
rect 115218 27922 115274 27978
rect 115342 27922 115398 27978
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 58294 129306 58350
rect 129374 58294 129430 58350
rect 129498 58294 129554 58350
rect 129622 58294 129678 58350
rect 129250 58170 129306 58226
rect 129374 58170 129430 58226
rect 129498 58170 129554 58226
rect 129622 58170 129678 58226
rect 129250 58046 129306 58102
rect 129374 58046 129430 58102
rect 129498 58046 129554 58102
rect 129622 58046 129678 58102
rect 129250 57922 129306 57978
rect 129374 57922 129430 57978
rect 129498 57922 129554 57978
rect 129622 57922 129678 57978
rect 129250 40294 129306 40350
rect 129374 40294 129430 40350
rect 129498 40294 129554 40350
rect 129622 40294 129678 40350
rect 129250 40170 129306 40226
rect 129374 40170 129430 40226
rect 129498 40170 129554 40226
rect 129622 40170 129678 40226
rect 129250 40046 129306 40102
rect 129374 40046 129430 40102
rect 129498 40046 129554 40102
rect 129622 40046 129678 40102
rect 129250 39922 129306 39978
rect 129374 39922 129430 39978
rect 129498 39922 129554 39978
rect 129622 39922 129678 39978
rect 129250 22294 129306 22350
rect 129374 22294 129430 22350
rect 129498 22294 129554 22350
rect 129622 22294 129678 22350
rect 129250 22170 129306 22226
rect 129374 22170 129430 22226
rect 129498 22170 129554 22226
rect 129622 22170 129678 22226
rect 129250 22046 129306 22102
rect 129374 22046 129430 22102
rect 129498 22046 129554 22102
rect 129622 22046 129678 22102
rect 129250 21922 129306 21978
rect 129374 21922 129430 21978
rect 129498 21922 129554 21978
rect 129622 21922 129678 21978
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 46294 133026 46350
rect 133094 46294 133150 46350
rect 133218 46294 133274 46350
rect 133342 46294 133398 46350
rect 132970 46170 133026 46226
rect 133094 46170 133150 46226
rect 133218 46170 133274 46226
rect 133342 46170 133398 46226
rect 132970 46046 133026 46102
rect 133094 46046 133150 46102
rect 133218 46046 133274 46102
rect 133342 46046 133398 46102
rect 132970 45922 133026 45978
rect 133094 45922 133150 45978
rect 133218 45922 133274 45978
rect 133342 45922 133398 45978
rect 132970 28294 133026 28350
rect 133094 28294 133150 28350
rect 133218 28294 133274 28350
rect 133342 28294 133398 28350
rect 132970 28170 133026 28226
rect 133094 28170 133150 28226
rect 133218 28170 133274 28226
rect 133342 28170 133398 28226
rect 132970 28046 133026 28102
rect 133094 28046 133150 28102
rect 133218 28046 133274 28102
rect 133342 28046 133398 28102
rect 132970 27922 133026 27978
rect 133094 27922 133150 27978
rect 133218 27922 133274 27978
rect 133342 27922 133398 27978
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 147250 58294 147306 58350
rect 147374 58294 147430 58350
rect 147498 58294 147554 58350
rect 147622 58294 147678 58350
rect 147250 58170 147306 58226
rect 147374 58170 147430 58226
rect 147498 58170 147554 58226
rect 147622 58170 147678 58226
rect 147250 58046 147306 58102
rect 147374 58046 147430 58102
rect 147498 58046 147554 58102
rect 147622 58046 147678 58102
rect 147250 57922 147306 57978
rect 147374 57922 147430 57978
rect 147498 57922 147554 57978
rect 147622 57922 147678 57978
rect 147250 40294 147306 40350
rect 147374 40294 147430 40350
rect 147498 40294 147554 40350
rect 147622 40294 147678 40350
rect 147250 40170 147306 40226
rect 147374 40170 147430 40226
rect 147498 40170 147554 40226
rect 147622 40170 147678 40226
rect 147250 40046 147306 40102
rect 147374 40046 147430 40102
rect 147498 40046 147554 40102
rect 147622 40046 147678 40102
rect 147250 39922 147306 39978
rect 147374 39922 147430 39978
rect 147498 39922 147554 39978
rect 147622 39922 147678 39978
rect 147250 22294 147306 22350
rect 147374 22294 147430 22350
rect 147498 22294 147554 22350
rect 147622 22294 147678 22350
rect 147250 22170 147306 22226
rect 147374 22170 147430 22226
rect 147498 22170 147554 22226
rect 147622 22170 147678 22226
rect 147250 22046 147306 22102
rect 147374 22046 147430 22102
rect 147498 22046 147554 22102
rect 147622 22046 147678 22102
rect 147250 21922 147306 21978
rect 147374 21922 147430 21978
rect 147498 21922 147554 21978
rect 147622 21922 147678 21978
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 150970 46294 151026 46350
rect 151094 46294 151150 46350
rect 151218 46294 151274 46350
rect 151342 46294 151398 46350
rect 150970 46170 151026 46226
rect 151094 46170 151150 46226
rect 151218 46170 151274 46226
rect 151342 46170 151398 46226
rect 150970 46046 151026 46102
rect 151094 46046 151150 46102
rect 151218 46046 151274 46102
rect 151342 46046 151398 46102
rect 150970 45922 151026 45978
rect 151094 45922 151150 45978
rect 151218 45922 151274 45978
rect 151342 45922 151398 45978
rect 150970 28294 151026 28350
rect 151094 28294 151150 28350
rect 151218 28294 151274 28350
rect 151342 28294 151398 28350
rect 150970 28170 151026 28226
rect 151094 28170 151150 28226
rect 151218 28170 151274 28226
rect 151342 28170 151398 28226
rect 150970 28046 151026 28102
rect 151094 28046 151150 28102
rect 151218 28046 151274 28102
rect 151342 28046 151398 28102
rect 150970 27922 151026 27978
rect 151094 27922 151150 27978
rect 151218 27922 151274 27978
rect 151342 27922 151398 27978
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 58294 165306 58350
rect 165374 58294 165430 58350
rect 165498 58294 165554 58350
rect 165622 58294 165678 58350
rect 165250 58170 165306 58226
rect 165374 58170 165430 58226
rect 165498 58170 165554 58226
rect 165622 58170 165678 58226
rect 165250 58046 165306 58102
rect 165374 58046 165430 58102
rect 165498 58046 165554 58102
rect 165622 58046 165678 58102
rect 165250 57922 165306 57978
rect 165374 57922 165430 57978
rect 165498 57922 165554 57978
rect 165622 57922 165678 57978
rect 165250 40294 165306 40350
rect 165374 40294 165430 40350
rect 165498 40294 165554 40350
rect 165622 40294 165678 40350
rect 165250 40170 165306 40226
rect 165374 40170 165430 40226
rect 165498 40170 165554 40226
rect 165622 40170 165678 40226
rect 165250 40046 165306 40102
rect 165374 40046 165430 40102
rect 165498 40046 165554 40102
rect 165622 40046 165678 40102
rect 165250 39922 165306 39978
rect 165374 39922 165430 39978
rect 165498 39922 165554 39978
rect 165622 39922 165678 39978
rect 165250 22294 165306 22350
rect 165374 22294 165430 22350
rect 165498 22294 165554 22350
rect 165622 22294 165678 22350
rect 165250 22170 165306 22226
rect 165374 22170 165430 22226
rect 165498 22170 165554 22226
rect 165622 22170 165678 22226
rect 165250 22046 165306 22102
rect 165374 22046 165430 22102
rect 165498 22046 165554 22102
rect 165622 22046 165678 22102
rect 165250 21922 165306 21978
rect 165374 21922 165430 21978
rect 165498 21922 165554 21978
rect 165622 21922 165678 21978
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 46294 169026 46350
rect 169094 46294 169150 46350
rect 169218 46294 169274 46350
rect 169342 46294 169398 46350
rect 168970 46170 169026 46226
rect 169094 46170 169150 46226
rect 169218 46170 169274 46226
rect 169342 46170 169398 46226
rect 168970 46046 169026 46102
rect 169094 46046 169150 46102
rect 169218 46046 169274 46102
rect 169342 46046 169398 46102
rect 168970 45922 169026 45978
rect 169094 45922 169150 45978
rect 169218 45922 169274 45978
rect 169342 45922 169398 45978
rect 168970 28294 169026 28350
rect 169094 28294 169150 28350
rect 169218 28294 169274 28350
rect 169342 28294 169398 28350
rect 168970 28170 169026 28226
rect 169094 28170 169150 28226
rect 169218 28170 169274 28226
rect 169342 28170 169398 28226
rect 168970 28046 169026 28102
rect 169094 28046 169150 28102
rect 169218 28046 169274 28102
rect 169342 28046 169398 28102
rect 168970 27922 169026 27978
rect 169094 27922 169150 27978
rect 169218 27922 169274 27978
rect 169342 27922 169398 27978
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 183250 58294 183306 58350
rect 183374 58294 183430 58350
rect 183498 58294 183554 58350
rect 183622 58294 183678 58350
rect 183250 58170 183306 58226
rect 183374 58170 183430 58226
rect 183498 58170 183554 58226
rect 183622 58170 183678 58226
rect 183250 58046 183306 58102
rect 183374 58046 183430 58102
rect 183498 58046 183554 58102
rect 183622 58046 183678 58102
rect 183250 57922 183306 57978
rect 183374 57922 183430 57978
rect 183498 57922 183554 57978
rect 183622 57922 183678 57978
rect 183250 40294 183306 40350
rect 183374 40294 183430 40350
rect 183498 40294 183554 40350
rect 183622 40294 183678 40350
rect 183250 40170 183306 40226
rect 183374 40170 183430 40226
rect 183498 40170 183554 40226
rect 183622 40170 183678 40226
rect 183250 40046 183306 40102
rect 183374 40046 183430 40102
rect 183498 40046 183554 40102
rect 183622 40046 183678 40102
rect 183250 39922 183306 39978
rect 183374 39922 183430 39978
rect 183498 39922 183554 39978
rect 183622 39922 183678 39978
rect 183250 22294 183306 22350
rect 183374 22294 183430 22350
rect 183498 22294 183554 22350
rect 183622 22294 183678 22350
rect 183250 22170 183306 22226
rect 183374 22170 183430 22226
rect 183498 22170 183554 22226
rect 183622 22170 183678 22226
rect 183250 22046 183306 22102
rect 183374 22046 183430 22102
rect 183498 22046 183554 22102
rect 183622 22046 183678 22102
rect 183250 21922 183306 21978
rect 183374 21922 183430 21978
rect 183498 21922 183554 21978
rect 183622 21922 183678 21978
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 46294 187026 46350
rect 187094 46294 187150 46350
rect 187218 46294 187274 46350
rect 187342 46294 187398 46350
rect 186970 46170 187026 46226
rect 187094 46170 187150 46226
rect 187218 46170 187274 46226
rect 187342 46170 187398 46226
rect 186970 46046 187026 46102
rect 187094 46046 187150 46102
rect 187218 46046 187274 46102
rect 187342 46046 187398 46102
rect 186970 45922 187026 45978
rect 187094 45922 187150 45978
rect 187218 45922 187274 45978
rect 187342 45922 187398 45978
rect 186970 28294 187026 28350
rect 187094 28294 187150 28350
rect 187218 28294 187274 28350
rect 187342 28294 187398 28350
rect 186970 28170 187026 28226
rect 187094 28170 187150 28226
rect 187218 28170 187274 28226
rect 187342 28170 187398 28226
rect 186970 28046 187026 28102
rect 187094 28046 187150 28102
rect 187218 28046 187274 28102
rect 187342 28046 187398 28102
rect 186970 27922 187026 27978
rect 187094 27922 187150 27978
rect 187218 27922 187274 27978
rect 187342 27922 187398 27978
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 201250 58294 201306 58350
rect 201374 58294 201430 58350
rect 201498 58294 201554 58350
rect 201622 58294 201678 58350
rect 201250 58170 201306 58226
rect 201374 58170 201430 58226
rect 201498 58170 201554 58226
rect 201622 58170 201678 58226
rect 201250 58046 201306 58102
rect 201374 58046 201430 58102
rect 201498 58046 201554 58102
rect 201622 58046 201678 58102
rect 201250 57922 201306 57978
rect 201374 57922 201430 57978
rect 201498 57922 201554 57978
rect 201622 57922 201678 57978
rect 201250 40294 201306 40350
rect 201374 40294 201430 40350
rect 201498 40294 201554 40350
rect 201622 40294 201678 40350
rect 201250 40170 201306 40226
rect 201374 40170 201430 40226
rect 201498 40170 201554 40226
rect 201622 40170 201678 40226
rect 201250 40046 201306 40102
rect 201374 40046 201430 40102
rect 201498 40046 201554 40102
rect 201622 40046 201678 40102
rect 201250 39922 201306 39978
rect 201374 39922 201430 39978
rect 201498 39922 201554 39978
rect 201622 39922 201678 39978
rect 201250 22294 201306 22350
rect 201374 22294 201430 22350
rect 201498 22294 201554 22350
rect 201622 22294 201678 22350
rect 201250 22170 201306 22226
rect 201374 22170 201430 22226
rect 201498 22170 201554 22226
rect 201622 22170 201678 22226
rect 201250 22046 201306 22102
rect 201374 22046 201430 22102
rect 201498 22046 201554 22102
rect 201622 22046 201678 22102
rect 201250 21922 201306 21978
rect 201374 21922 201430 21978
rect 201498 21922 201554 21978
rect 201622 21922 201678 21978
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 204970 46294 205026 46350
rect 205094 46294 205150 46350
rect 205218 46294 205274 46350
rect 205342 46294 205398 46350
rect 204970 46170 205026 46226
rect 205094 46170 205150 46226
rect 205218 46170 205274 46226
rect 205342 46170 205398 46226
rect 204970 46046 205026 46102
rect 205094 46046 205150 46102
rect 205218 46046 205274 46102
rect 205342 46046 205398 46102
rect 204970 45922 205026 45978
rect 205094 45922 205150 45978
rect 205218 45922 205274 45978
rect 205342 45922 205398 45978
rect 204970 28294 205026 28350
rect 205094 28294 205150 28350
rect 205218 28294 205274 28350
rect 205342 28294 205398 28350
rect 204970 28170 205026 28226
rect 205094 28170 205150 28226
rect 205218 28170 205274 28226
rect 205342 28170 205398 28226
rect 204970 28046 205026 28102
rect 205094 28046 205150 28102
rect 205218 28046 205274 28102
rect 205342 28046 205398 28102
rect 204970 27922 205026 27978
rect 205094 27922 205150 27978
rect 205218 27922 205274 27978
rect 205342 27922 205398 27978
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 219250 58294 219306 58350
rect 219374 58294 219430 58350
rect 219498 58294 219554 58350
rect 219622 58294 219678 58350
rect 219250 58170 219306 58226
rect 219374 58170 219430 58226
rect 219498 58170 219554 58226
rect 219622 58170 219678 58226
rect 219250 58046 219306 58102
rect 219374 58046 219430 58102
rect 219498 58046 219554 58102
rect 219622 58046 219678 58102
rect 219250 57922 219306 57978
rect 219374 57922 219430 57978
rect 219498 57922 219554 57978
rect 219622 57922 219678 57978
rect 219250 40294 219306 40350
rect 219374 40294 219430 40350
rect 219498 40294 219554 40350
rect 219622 40294 219678 40350
rect 219250 40170 219306 40226
rect 219374 40170 219430 40226
rect 219498 40170 219554 40226
rect 219622 40170 219678 40226
rect 219250 40046 219306 40102
rect 219374 40046 219430 40102
rect 219498 40046 219554 40102
rect 219622 40046 219678 40102
rect 219250 39922 219306 39978
rect 219374 39922 219430 39978
rect 219498 39922 219554 39978
rect 219622 39922 219678 39978
rect 219250 22294 219306 22350
rect 219374 22294 219430 22350
rect 219498 22294 219554 22350
rect 219622 22294 219678 22350
rect 219250 22170 219306 22226
rect 219374 22170 219430 22226
rect 219498 22170 219554 22226
rect 219622 22170 219678 22226
rect 219250 22046 219306 22102
rect 219374 22046 219430 22102
rect 219498 22046 219554 22102
rect 219622 22046 219678 22102
rect 219250 21922 219306 21978
rect 219374 21922 219430 21978
rect 219498 21922 219554 21978
rect 219622 21922 219678 21978
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 222970 46294 223026 46350
rect 223094 46294 223150 46350
rect 223218 46294 223274 46350
rect 223342 46294 223398 46350
rect 222970 46170 223026 46226
rect 223094 46170 223150 46226
rect 223218 46170 223274 46226
rect 223342 46170 223398 46226
rect 222970 46046 223026 46102
rect 223094 46046 223150 46102
rect 223218 46046 223274 46102
rect 223342 46046 223398 46102
rect 222970 45922 223026 45978
rect 223094 45922 223150 45978
rect 223218 45922 223274 45978
rect 223342 45922 223398 45978
rect 222970 28294 223026 28350
rect 223094 28294 223150 28350
rect 223218 28294 223274 28350
rect 223342 28294 223398 28350
rect 222970 28170 223026 28226
rect 223094 28170 223150 28226
rect 223218 28170 223274 28226
rect 223342 28170 223398 28226
rect 222970 28046 223026 28102
rect 223094 28046 223150 28102
rect 223218 28046 223274 28102
rect 223342 28046 223398 28102
rect 222970 27922 223026 27978
rect 223094 27922 223150 27978
rect 223218 27922 223274 27978
rect 223342 27922 223398 27978
rect 222970 10294 223026 10350
rect 223094 10294 223150 10350
rect 223218 10294 223274 10350
rect 223342 10294 223398 10350
rect 222970 10170 223026 10226
rect 223094 10170 223150 10226
rect 223218 10170 223274 10226
rect 223342 10170 223398 10226
rect 222970 10046 223026 10102
rect 223094 10046 223150 10102
rect 223218 10046 223274 10102
rect 223342 10046 223398 10102
rect 222970 9922 223026 9978
rect 223094 9922 223150 9978
rect 223218 9922 223274 9978
rect 223342 9922 223398 9978
rect 222970 -1176 223026 -1120
rect 223094 -1176 223150 -1120
rect 223218 -1176 223274 -1120
rect 223342 -1176 223398 -1120
rect 222970 -1300 223026 -1244
rect 223094 -1300 223150 -1244
rect 223218 -1300 223274 -1244
rect 223342 -1300 223398 -1244
rect 222970 -1424 223026 -1368
rect 223094 -1424 223150 -1368
rect 223218 -1424 223274 -1368
rect 223342 -1424 223398 -1368
rect 222970 -1548 223026 -1492
rect 223094 -1548 223150 -1492
rect 223218 -1548 223274 -1492
rect 223342 -1548 223398 -1492
rect 237250 58294 237306 58350
rect 237374 58294 237430 58350
rect 237498 58294 237554 58350
rect 237622 58294 237678 58350
rect 237250 58170 237306 58226
rect 237374 58170 237430 58226
rect 237498 58170 237554 58226
rect 237622 58170 237678 58226
rect 237250 58046 237306 58102
rect 237374 58046 237430 58102
rect 237498 58046 237554 58102
rect 237622 58046 237678 58102
rect 237250 57922 237306 57978
rect 237374 57922 237430 57978
rect 237498 57922 237554 57978
rect 237622 57922 237678 57978
rect 237250 40294 237306 40350
rect 237374 40294 237430 40350
rect 237498 40294 237554 40350
rect 237622 40294 237678 40350
rect 237250 40170 237306 40226
rect 237374 40170 237430 40226
rect 237498 40170 237554 40226
rect 237622 40170 237678 40226
rect 237250 40046 237306 40102
rect 237374 40046 237430 40102
rect 237498 40046 237554 40102
rect 237622 40046 237678 40102
rect 237250 39922 237306 39978
rect 237374 39922 237430 39978
rect 237498 39922 237554 39978
rect 237622 39922 237678 39978
rect 237250 22294 237306 22350
rect 237374 22294 237430 22350
rect 237498 22294 237554 22350
rect 237622 22294 237678 22350
rect 237250 22170 237306 22226
rect 237374 22170 237430 22226
rect 237498 22170 237554 22226
rect 237622 22170 237678 22226
rect 237250 22046 237306 22102
rect 237374 22046 237430 22102
rect 237498 22046 237554 22102
rect 237622 22046 237678 22102
rect 237250 21922 237306 21978
rect 237374 21922 237430 21978
rect 237498 21922 237554 21978
rect 237622 21922 237678 21978
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 240970 46294 241026 46350
rect 241094 46294 241150 46350
rect 241218 46294 241274 46350
rect 241342 46294 241398 46350
rect 240970 46170 241026 46226
rect 241094 46170 241150 46226
rect 241218 46170 241274 46226
rect 241342 46170 241398 46226
rect 240970 46046 241026 46102
rect 241094 46046 241150 46102
rect 241218 46046 241274 46102
rect 241342 46046 241398 46102
rect 240970 45922 241026 45978
rect 241094 45922 241150 45978
rect 241218 45922 241274 45978
rect 241342 45922 241398 45978
rect 240970 28294 241026 28350
rect 241094 28294 241150 28350
rect 241218 28294 241274 28350
rect 241342 28294 241398 28350
rect 240970 28170 241026 28226
rect 241094 28170 241150 28226
rect 241218 28170 241274 28226
rect 241342 28170 241398 28226
rect 240970 28046 241026 28102
rect 241094 28046 241150 28102
rect 241218 28046 241274 28102
rect 241342 28046 241398 28102
rect 240970 27922 241026 27978
rect 241094 27922 241150 27978
rect 241218 27922 241274 27978
rect 241342 27922 241398 27978
rect 240970 10294 241026 10350
rect 241094 10294 241150 10350
rect 241218 10294 241274 10350
rect 241342 10294 241398 10350
rect 240970 10170 241026 10226
rect 241094 10170 241150 10226
rect 241218 10170 241274 10226
rect 241342 10170 241398 10226
rect 240970 10046 241026 10102
rect 241094 10046 241150 10102
rect 241218 10046 241274 10102
rect 241342 10046 241398 10102
rect 240970 9922 241026 9978
rect 241094 9922 241150 9978
rect 241218 9922 241274 9978
rect 241342 9922 241398 9978
rect 240970 -1176 241026 -1120
rect 241094 -1176 241150 -1120
rect 241218 -1176 241274 -1120
rect 241342 -1176 241398 -1120
rect 240970 -1300 241026 -1244
rect 241094 -1300 241150 -1244
rect 241218 -1300 241274 -1244
rect 241342 -1300 241398 -1244
rect 240970 -1424 241026 -1368
rect 241094 -1424 241150 -1368
rect 241218 -1424 241274 -1368
rect 241342 -1424 241398 -1368
rect 240970 -1548 241026 -1492
rect 241094 -1548 241150 -1492
rect 241218 -1548 241274 -1492
rect 241342 -1548 241398 -1492
rect 255250 58294 255306 58350
rect 255374 58294 255430 58350
rect 255498 58294 255554 58350
rect 255622 58294 255678 58350
rect 255250 58170 255306 58226
rect 255374 58170 255430 58226
rect 255498 58170 255554 58226
rect 255622 58170 255678 58226
rect 255250 58046 255306 58102
rect 255374 58046 255430 58102
rect 255498 58046 255554 58102
rect 255622 58046 255678 58102
rect 255250 57922 255306 57978
rect 255374 57922 255430 57978
rect 255498 57922 255554 57978
rect 255622 57922 255678 57978
rect 255250 40294 255306 40350
rect 255374 40294 255430 40350
rect 255498 40294 255554 40350
rect 255622 40294 255678 40350
rect 255250 40170 255306 40226
rect 255374 40170 255430 40226
rect 255498 40170 255554 40226
rect 255622 40170 255678 40226
rect 255250 40046 255306 40102
rect 255374 40046 255430 40102
rect 255498 40046 255554 40102
rect 255622 40046 255678 40102
rect 255250 39922 255306 39978
rect 255374 39922 255430 39978
rect 255498 39922 255554 39978
rect 255622 39922 255678 39978
rect 255250 22294 255306 22350
rect 255374 22294 255430 22350
rect 255498 22294 255554 22350
rect 255622 22294 255678 22350
rect 255250 22170 255306 22226
rect 255374 22170 255430 22226
rect 255498 22170 255554 22226
rect 255622 22170 255678 22226
rect 255250 22046 255306 22102
rect 255374 22046 255430 22102
rect 255498 22046 255554 22102
rect 255622 22046 255678 22102
rect 255250 21922 255306 21978
rect 255374 21922 255430 21978
rect 255498 21922 255554 21978
rect 255622 21922 255678 21978
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 258970 46294 259026 46350
rect 259094 46294 259150 46350
rect 259218 46294 259274 46350
rect 259342 46294 259398 46350
rect 258970 46170 259026 46226
rect 259094 46170 259150 46226
rect 259218 46170 259274 46226
rect 259342 46170 259398 46226
rect 258970 46046 259026 46102
rect 259094 46046 259150 46102
rect 259218 46046 259274 46102
rect 259342 46046 259398 46102
rect 258970 45922 259026 45978
rect 259094 45922 259150 45978
rect 259218 45922 259274 45978
rect 259342 45922 259398 45978
rect 258970 28294 259026 28350
rect 259094 28294 259150 28350
rect 259218 28294 259274 28350
rect 259342 28294 259398 28350
rect 258970 28170 259026 28226
rect 259094 28170 259150 28226
rect 259218 28170 259274 28226
rect 259342 28170 259398 28226
rect 258970 28046 259026 28102
rect 259094 28046 259150 28102
rect 259218 28046 259274 28102
rect 259342 28046 259398 28102
rect 258970 27922 259026 27978
rect 259094 27922 259150 27978
rect 259218 27922 259274 27978
rect 259342 27922 259398 27978
rect 258970 10294 259026 10350
rect 259094 10294 259150 10350
rect 259218 10294 259274 10350
rect 259342 10294 259398 10350
rect 258970 10170 259026 10226
rect 259094 10170 259150 10226
rect 259218 10170 259274 10226
rect 259342 10170 259398 10226
rect 258970 10046 259026 10102
rect 259094 10046 259150 10102
rect 259218 10046 259274 10102
rect 259342 10046 259398 10102
rect 258970 9922 259026 9978
rect 259094 9922 259150 9978
rect 259218 9922 259274 9978
rect 259342 9922 259398 9978
rect 258970 -1176 259026 -1120
rect 259094 -1176 259150 -1120
rect 259218 -1176 259274 -1120
rect 259342 -1176 259398 -1120
rect 258970 -1300 259026 -1244
rect 259094 -1300 259150 -1244
rect 259218 -1300 259274 -1244
rect 259342 -1300 259398 -1244
rect 258970 -1424 259026 -1368
rect 259094 -1424 259150 -1368
rect 259218 -1424 259274 -1368
rect 259342 -1424 259398 -1368
rect 258970 -1548 259026 -1492
rect 259094 -1548 259150 -1492
rect 259218 -1548 259274 -1492
rect 259342 -1548 259398 -1492
rect 273250 58294 273306 58350
rect 273374 58294 273430 58350
rect 273498 58294 273554 58350
rect 273622 58294 273678 58350
rect 273250 58170 273306 58226
rect 273374 58170 273430 58226
rect 273498 58170 273554 58226
rect 273622 58170 273678 58226
rect 273250 58046 273306 58102
rect 273374 58046 273430 58102
rect 273498 58046 273554 58102
rect 273622 58046 273678 58102
rect 273250 57922 273306 57978
rect 273374 57922 273430 57978
rect 273498 57922 273554 57978
rect 273622 57922 273678 57978
rect 273250 40294 273306 40350
rect 273374 40294 273430 40350
rect 273498 40294 273554 40350
rect 273622 40294 273678 40350
rect 273250 40170 273306 40226
rect 273374 40170 273430 40226
rect 273498 40170 273554 40226
rect 273622 40170 273678 40226
rect 273250 40046 273306 40102
rect 273374 40046 273430 40102
rect 273498 40046 273554 40102
rect 273622 40046 273678 40102
rect 273250 39922 273306 39978
rect 273374 39922 273430 39978
rect 273498 39922 273554 39978
rect 273622 39922 273678 39978
rect 273250 22294 273306 22350
rect 273374 22294 273430 22350
rect 273498 22294 273554 22350
rect 273622 22294 273678 22350
rect 273250 22170 273306 22226
rect 273374 22170 273430 22226
rect 273498 22170 273554 22226
rect 273622 22170 273678 22226
rect 273250 22046 273306 22102
rect 273374 22046 273430 22102
rect 273498 22046 273554 22102
rect 273622 22046 273678 22102
rect 273250 21922 273306 21978
rect 273374 21922 273430 21978
rect 273498 21922 273554 21978
rect 273622 21922 273678 21978
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 276970 46294 277026 46350
rect 277094 46294 277150 46350
rect 277218 46294 277274 46350
rect 277342 46294 277398 46350
rect 276970 46170 277026 46226
rect 277094 46170 277150 46226
rect 277218 46170 277274 46226
rect 277342 46170 277398 46226
rect 276970 46046 277026 46102
rect 277094 46046 277150 46102
rect 277218 46046 277274 46102
rect 277342 46046 277398 46102
rect 276970 45922 277026 45978
rect 277094 45922 277150 45978
rect 277218 45922 277274 45978
rect 277342 45922 277398 45978
rect 276970 28294 277026 28350
rect 277094 28294 277150 28350
rect 277218 28294 277274 28350
rect 277342 28294 277398 28350
rect 276970 28170 277026 28226
rect 277094 28170 277150 28226
rect 277218 28170 277274 28226
rect 277342 28170 277398 28226
rect 276970 28046 277026 28102
rect 277094 28046 277150 28102
rect 277218 28046 277274 28102
rect 277342 28046 277398 28102
rect 276970 27922 277026 27978
rect 277094 27922 277150 27978
rect 277218 27922 277274 27978
rect 277342 27922 277398 27978
rect 276970 10294 277026 10350
rect 277094 10294 277150 10350
rect 277218 10294 277274 10350
rect 277342 10294 277398 10350
rect 276970 10170 277026 10226
rect 277094 10170 277150 10226
rect 277218 10170 277274 10226
rect 277342 10170 277398 10226
rect 276970 10046 277026 10102
rect 277094 10046 277150 10102
rect 277218 10046 277274 10102
rect 277342 10046 277398 10102
rect 276970 9922 277026 9978
rect 277094 9922 277150 9978
rect 277218 9922 277274 9978
rect 277342 9922 277398 9978
rect 276970 -1176 277026 -1120
rect 277094 -1176 277150 -1120
rect 277218 -1176 277274 -1120
rect 277342 -1176 277398 -1120
rect 276970 -1300 277026 -1244
rect 277094 -1300 277150 -1244
rect 277218 -1300 277274 -1244
rect 277342 -1300 277398 -1244
rect 276970 -1424 277026 -1368
rect 277094 -1424 277150 -1368
rect 277218 -1424 277274 -1368
rect 277342 -1424 277398 -1368
rect 276970 -1548 277026 -1492
rect 277094 -1548 277150 -1492
rect 277218 -1548 277274 -1492
rect 277342 -1548 277398 -1492
rect 291250 58294 291306 58350
rect 291374 58294 291430 58350
rect 291498 58294 291554 58350
rect 291622 58294 291678 58350
rect 291250 58170 291306 58226
rect 291374 58170 291430 58226
rect 291498 58170 291554 58226
rect 291622 58170 291678 58226
rect 291250 58046 291306 58102
rect 291374 58046 291430 58102
rect 291498 58046 291554 58102
rect 291622 58046 291678 58102
rect 291250 57922 291306 57978
rect 291374 57922 291430 57978
rect 291498 57922 291554 57978
rect 291622 57922 291678 57978
rect 291250 40294 291306 40350
rect 291374 40294 291430 40350
rect 291498 40294 291554 40350
rect 291622 40294 291678 40350
rect 291250 40170 291306 40226
rect 291374 40170 291430 40226
rect 291498 40170 291554 40226
rect 291622 40170 291678 40226
rect 291250 40046 291306 40102
rect 291374 40046 291430 40102
rect 291498 40046 291554 40102
rect 291622 40046 291678 40102
rect 291250 39922 291306 39978
rect 291374 39922 291430 39978
rect 291498 39922 291554 39978
rect 291622 39922 291678 39978
rect 291250 22294 291306 22350
rect 291374 22294 291430 22350
rect 291498 22294 291554 22350
rect 291622 22294 291678 22350
rect 291250 22170 291306 22226
rect 291374 22170 291430 22226
rect 291498 22170 291554 22226
rect 291622 22170 291678 22226
rect 291250 22046 291306 22102
rect 291374 22046 291430 22102
rect 291498 22046 291554 22102
rect 291622 22046 291678 22102
rect 291250 21922 291306 21978
rect 291374 21922 291430 21978
rect 291498 21922 291554 21978
rect 291622 21922 291678 21978
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 294970 46294 295026 46350
rect 295094 46294 295150 46350
rect 295218 46294 295274 46350
rect 295342 46294 295398 46350
rect 294970 46170 295026 46226
rect 295094 46170 295150 46226
rect 295218 46170 295274 46226
rect 295342 46170 295398 46226
rect 294970 46046 295026 46102
rect 295094 46046 295150 46102
rect 295218 46046 295274 46102
rect 295342 46046 295398 46102
rect 294970 45922 295026 45978
rect 295094 45922 295150 45978
rect 295218 45922 295274 45978
rect 295342 45922 295398 45978
rect 294970 28294 295026 28350
rect 295094 28294 295150 28350
rect 295218 28294 295274 28350
rect 295342 28294 295398 28350
rect 294970 28170 295026 28226
rect 295094 28170 295150 28226
rect 295218 28170 295274 28226
rect 295342 28170 295398 28226
rect 294970 28046 295026 28102
rect 295094 28046 295150 28102
rect 295218 28046 295274 28102
rect 295342 28046 295398 28102
rect 294970 27922 295026 27978
rect 295094 27922 295150 27978
rect 295218 27922 295274 27978
rect 295342 27922 295398 27978
rect 294970 10294 295026 10350
rect 295094 10294 295150 10350
rect 295218 10294 295274 10350
rect 295342 10294 295398 10350
rect 294970 10170 295026 10226
rect 295094 10170 295150 10226
rect 295218 10170 295274 10226
rect 295342 10170 295398 10226
rect 294970 10046 295026 10102
rect 295094 10046 295150 10102
rect 295218 10046 295274 10102
rect 295342 10046 295398 10102
rect 294970 9922 295026 9978
rect 295094 9922 295150 9978
rect 295218 9922 295274 9978
rect 295342 9922 295398 9978
rect 294970 -1176 295026 -1120
rect 295094 -1176 295150 -1120
rect 295218 -1176 295274 -1120
rect 295342 -1176 295398 -1120
rect 294970 -1300 295026 -1244
rect 295094 -1300 295150 -1244
rect 295218 -1300 295274 -1244
rect 295342 -1300 295398 -1244
rect 294970 -1424 295026 -1368
rect 295094 -1424 295150 -1368
rect 295218 -1424 295274 -1368
rect 295342 -1424 295398 -1368
rect 294970 -1548 295026 -1492
rect 295094 -1548 295150 -1492
rect 295218 -1548 295274 -1492
rect 295342 -1548 295398 -1492
rect 309250 58294 309306 58350
rect 309374 58294 309430 58350
rect 309498 58294 309554 58350
rect 309622 58294 309678 58350
rect 309250 58170 309306 58226
rect 309374 58170 309430 58226
rect 309498 58170 309554 58226
rect 309622 58170 309678 58226
rect 309250 58046 309306 58102
rect 309374 58046 309430 58102
rect 309498 58046 309554 58102
rect 309622 58046 309678 58102
rect 309250 57922 309306 57978
rect 309374 57922 309430 57978
rect 309498 57922 309554 57978
rect 309622 57922 309678 57978
rect 309250 40294 309306 40350
rect 309374 40294 309430 40350
rect 309498 40294 309554 40350
rect 309622 40294 309678 40350
rect 309250 40170 309306 40226
rect 309374 40170 309430 40226
rect 309498 40170 309554 40226
rect 309622 40170 309678 40226
rect 309250 40046 309306 40102
rect 309374 40046 309430 40102
rect 309498 40046 309554 40102
rect 309622 40046 309678 40102
rect 309250 39922 309306 39978
rect 309374 39922 309430 39978
rect 309498 39922 309554 39978
rect 309622 39922 309678 39978
rect 309250 22294 309306 22350
rect 309374 22294 309430 22350
rect 309498 22294 309554 22350
rect 309622 22294 309678 22350
rect 309250 22170 309306 22226
rect 309374 22170 309430 22226
rect 309498 22170 309554 22226
rect 309622 22170 309678 22226
rect 309250 22046 309306 22102
rect 309374 22046 309430 22102
rect 309498 22046 309554 22102
rect 309622 22046 309678 22102
rect 309250 21922 309306 21978
rect 309374 21922 309430 21978
rect 309498 21922 309554 21978
rect 309622 21922 309678 21978
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 312970 46294 313026 46350
rect 313094 46294 313150 46350
rect 313218 46294 313274 46350
rect 313342 46294 313398 46350
rect 312970 46170 313026 46226
rect 313094 46170 313150 46226
rect 313218 46170 313274 46226
rect 313342 46170 313398 46226
rect 312970 46046 313026 46102
rect 313094 46046 313150 46102
rect 313218 46046 313274 46102
rect 313342 46046 313398 46102
rect 312970 45922 313026 45978
rect 313094 45922 313150 45978
rect 313218 45922 313274 45978
rect 313342 45922 313398 45978
rect 312970 28294 313026 28350
rect 313094 28294 313150 28350
rect 313218 28294 313274 28350
rect 313342 28294 313398 28350
rect 312970 28170 313026 28226
rect 313094 28170 313150 28226
rect 313218 28170 313274 28226
rect 313342 28170 313398 28226
rect 312970 28046 313026 28102
rect 313094 28046 313150 28102
rect 313218 28046 313274 28102
rect 313342 28046 313398 28102
rect 312970 27922 313026 27978
rect 313094 27922 313150 27978
rect 313218 27922 313274 27978
rect 313342 27922 313398 27978
rect 312970 10294 313026 10350
rect 313094 10294 313150 10350
rect 313218 10294 313274 10350
rect 313342 10294 313398 10350
rect 312970 10170 313026 10226
rect 313094 10170 313150 10226
rect 313218 10170 313274 10226
rect 313342 10170 313398 10226
rect 312970 10046 313026 10102
rect 313094 10046 313150 10102
rect 313218 10046 313274 10102
rect 313342 10046 313398 10102
rect 312970 9922 313026 9978
rect 313094 9922 313150 9978
rect 313218 9922 313274 9978
rect 313342 9922 313398 9978
rect 312970 -1176 313026 -1120
rect 313094 -1176 313150 -1120
rect 313218 -1176 313274 -1120
rect 313342 -1176 313398 -1120
rect 312970 -1300 313026 -1244
rect 313094 -1300 313150 -1244
rect 313218 -1300 313274 -1244
rect 313342 -1300 313398 -1244
rect 312970 -1424 313026 -1368
rect 313094 -1424 313150 -1368
rect 313218 -1424 313274 -1368
rect 313342 -1424 313398 -1368
rect 312970 -1548 313026 -1492
rect 313094 -1548 313150 -1492
rect 313218 -1548 313274 -1492
rect 313342 -1548 313398 -1492
rect 327250 58294 327306 58350
rect 327374 58294 327430 58350
rect 327498 58294 327554 58350
rect 327622 58294 327678 58350
rect 327250 58170 327306 58226
rect 327374 58170 327430 58226
rect 327498 58170 327554 58226
rect 327622 58170 327678 58226
rect 327250 58046 327306 58102
rect 327374 58046 327430 58102
rect 327498 58046 327554 58102
rect 327622 58046 327678 58102
rect 327250 57922 327306 57978
rect 327374 57922 327430 57978
rect 327498 57922 327554 57978
rect 327622 57922 327678 57978
rect 327250 40294 327306 40350
rect 327374 40294 327430 40350
rect 327498 40294 327554 40350
rect 327622 40294 327678 40350
rect 327250 40170 327306 40226
rect 327374 40170 327430 40226
rect 327498 40170 327554 40226
rect 327622 40170 327678 40226
rect 327250 40046 327306 40102
rect 327374 40046 327430 40102
rect 327498 40046 327554 40102
rect 327622 40046 327678 40102
rect 327250 39922 327306 39978
rect 327374 39922 327430 39978
rect 327498 39922 327554 39978
rect 327622 39922 327678 39978
rect 327250 22294 327306 22350
rect 327374 22294 327430 22350
rect 327498 22294 327554 22350
rect 327622 22294 327678 22350
rect 327250 22170 327306 22226
rect 327374 22170 327430 22226
rect 327498 22170 327554 22226
rect 327622 22170 327678 22226
rect 327250 22046 327306 22102
rect 327374 22046 327430 22102
rect 327498 22046 327554 22102
rect 327622 22046 327678 22102
rect 327250 21922 327306 21978
rect 327374 21922 327430 21978
rect 327498 21922 327554 21978
rect 327622 21922 327678 21978
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 330970 46294 331026 46350
rect 331094 46294 331150 46350
rect 331218 46294 331274 46350
rect 331342 46294 331398 46350
rect 330970 46170 331026 46226
rect 331094 46170 331150 46226
rect 331218 46170 331274 46226
rect 331342 46170 331398 46226
rect 330970 46046 331026 46102
rect 331094 46046 331150 46102
rect 331218 46046 331274 46102
rect 331342 46046 331398 46102
rect 330970 45922 331026 45978
rect 331094 45922 331150 45978
rect 331218 45922 331274 45978
rect 331342 45922 331398 45978
rect 330970 28294 331026 28350
rect 331094 28294 331150 28350
rect 331218 28294 331274 28350
rect 331342 28294 331398 28350
rect 330970 28170 331026 28226
rect 331094 28170 331150 28226
rect 331218 28170 331274 28226
rect 331342 28170 331398 28226
rect 330970 28046 331026 28102
rect 331094 28046 331150 28102
rect 331218 28046 331274 28102
rect 331342 28046 331398 28102
rect 330970 27922 331026 27978
rect 331094 27922 331150 27978
rect 331218 27922 331274 27978
rect 331342 27922 331398 27978
rect 330970 10294 331026 10350
rect 331094 10294 331150 10350
rect 331218 10294 331274 10350
rect 331342 10294 331398 10350
rect 330970 10170 331026 10226
rect 331094 10170 331150 10226
rect 331218 10170 331274 10226
rect 331342 10170 331398 10226
rect 330970 10046 331026 10102
rect 331094 10046 331150 10102
rect 331218 10046 331274 10102
rect 331342 10046 331398 10102
rect 330970 9922 331026 9978
rect 331094 9922 331150 9978
rect 331218 9922 331274 9978
rect 331342 9922 331398 9978
rect 330970 -1176 331026 -1120
rect 331094 -1176 331150 -1120
rect 331218 -1176 331274 -1120
rect 331342 -1176 331398 -1120
rect 330970 -1300 331026 -1244
rect 331094 -1300 331150 -1244
rect 331218 -1300 331274 -1244
rect 331342 -1300 331398 -1244
rect 330970 -1424 331026 -1368
rect 331094 -1424 331150 -1368
rect 331218 -1424 331274 -1368
rect 331342 -1424 331398 -1368
rect 330970 -1548 331026 -1492
rect 331094 -1548 331150 -1492
rect 331218 -1548 331274 -1492
rect 331342 -1548 331398 -1492
rect 345250 58294 345306 58350
rect 345374 58294 345430 58350
rect 345498 58294 345554 58350
rect 345622 58294 345678 58350
rect 345250 58170 345306 58226
rect 345374 58170 345430 58226
rect 345498 58170 345554 58226
rect 345622 58170 345678 58226
rect 345250 58046 345306 58102
rect 345374 58046 345430 58102
rect 345498 58046 345554 58102
rect 345622 58046 345678 58102
rect 345250 57922 345306 57978
rect 345374 57922 345430 57978
rect 345498 57922 345554 57978
rect 345622 57922 345678 57978
rect 345250 40294 345306 40350
rect 345374 40294 345430 40350
rect 345498 40294 345554 40350
rect 345622 40294 345678 40350
rect 345250 40170 345306 40226
rect 345374 40170 345430 40226
rect 345498 40170 345554 40226
rect 345622 40170 345678 40226
rect 345250 40046 345306 40102
rect 345374 40046 345430 40102
rect 345498 40046 345554 40102
rect 345622 40046 345678 40102
rect 345250 39922 345306 39978
rect 345374 39922 345430 39978
rect 345498 39922 345554 39978
rect 345622 39922 345678 39978
rect 345250 22294 345306 22350
rect 345374 22294 345430 22350
rect 345498 22294 345554 22350
rect 345622 22294 345678 22350
rect 345250 22170 345306 22226
rect 345374 22170 345430 22226
rect 345498 22170 345554 22226
rect 345622 22170 345678 22226
rect 345250 22046 345306 22102
rect 345374 22046 345430 22102
rect 345498 22046 345554 22102
rect 345622 22046 345678 22102
rect 345250 21922 345306 21978
rect 345374 21922 345430 21978
rect 345498 21922 345554 21978
rect 345622 21922 345678 21978
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 356358 64294 356414 64350
rect 356482 64294 356538 64350
rect 356358 64170 356414 64226
rect 356482 64170 356538 64226
rect 356358 64046 356414 64102
rect 356482 64046 356538 64102
rect 356358 63922 356414 63978
rect 356482 63922 356538 63978
rect 348970 46294 349026 46350
rect 349094 46294 349150 46350
rect 349218 46294 349274 46350
rect 349342 46294 349398 46350
rect 348970 46170 349026 46226
rect 349094 46170 349150 46226
rect 349218 46170 349274 46226
rect 349342 46170 349398 46226
rect 348970 46046 349026 46102
rect 349094 46046 349150 46102
rect 349218 46046 349274 46102
rect 349342 46046 349398 46102
rect 348970 45922 349026 45978
rect 349094 45922 349150 45978
rect 349218 45922 349274 45978
rect 349342 45922 349398 45978
rect 348970 28294 349026 28350
rect 349094 28294 349150 28350
rect 349218 28294 349274 28350
rect 349342 28294 349398 28350
rect 348970 28170 349026 28226
rect 349094 28170 349150 28226
rect 349218 28170 349274 28226
rect 349342 28170 349398 28226
rect 348970 28046 349026 28102
rect 349094 28046 349150 28102
rect 349218 28046 349274 28102
rect 349342 28046 349398 28102
rect 348970 27922 349026 27978
rect 349094 27922 349150 27978
rect 349218 27922 349274 27978
rect 349342 27922 349398 27978
rect 348970 10294 349026 10350
rect 349094 10294 349150 10350
rect 349218 10294 349274 10350
rect 349342 10294 349398 10350
rect 348970 10170 349026 10226
rect 349094 10170 349150 10226
rect 349218 10170 349274 10226
rect 349342 10170 349398 10226
rect 348970 10046 349026 10102
rect 349094 10046 349150 10102
rect 349218 10046 349274 10102
rect 349342 10046 349398 10102
rect 348970 9922 349026 9978
rect 349094 9922 349150 9978
rect 349218 9922 349274 9978
rect 349342 9922 349398 9978
rect 348970 -1176 349026 -1120
rect 349094 -1176 349150 -1120
rect 349218 -1176 349274 -1120
rect 349342 -1176 349398 -1120
rect 348970 -1300 349026 -1244
rect 349094 -1300 349150 -1244
rect 349218 -1300 349274 -1244
rect 349342 -1300 349398 -1244
rect 348970 -1424 349026 -1368
rect 349094 -1424 349150 -1368
rect 349218 -1424 349274 -1368
rect 349342 -1424 349398 -1368
rect 348970 -1548 349026 -1492
rect 349094 -1548 349150 -1492
rect 349218 -1548 349274 -1492
rect 349342 -1548 349398 -1492
rect 363250 58294 363306 58350
rect 363374 58294 363430 58350
rect 363498 58294 363554 58350
rect 363622 58294 363678 58350
rect 363250 58170 363306 58226
rect 363374 58170 363430 58226
rect 363498 58170 363554 58226
rect 363622 58170 363678 58226
rect 363250 58046 363306 58102
rect 363374 58046 363430 58102
rect 363498 58046 363554 58102
rect 363622 58046 363678 58102
rect 363250 57922 363306 57978
rect 363374 57922 363430 57978
rect 363498 57922 363554 57978
rect 363622 57922 363678 57978
rect 363250 40294 363306 40350
rect 363374 40294 363430 40350
rect 363498 40294 363554 40350
rect 363622 40294 363678 40350
rect 363250 40170 363306 40226
rect 363374 40170 363430 40226
rect 363498 40170 363554 40226
rect 363622 40170 363678 40226
rect 363250 40046 363306 40102
rect 363374 40046 363430 40102
rect 363498 40046 363554 40102
rect 363622 40046 363678 40102
rect 363250 39922 363306 39978
rect 363374 39922 363430 39978
rect 363498 39922 363554 39978
rect 363622 39922 363678 39978
rect 363250 22294 363306 22350
rect 363374 22294 363430 22350
rect 363498 22294 363554 22350
rect 363622 22294 363678 22350
rect 363250 22170 363306 22226
rect 363374 22170 363430 22226
rect 363498 22170 363554 22226
rect 363622 22170 363678 22226
rect 363250 22046 363306 22102
rect 363374 22046 363430 22102
rect 363498 22046 363554 22102
rect 363622 22046 363678 22102
rect 363250 21922 363306 21978
rect 363374 21922 363430 21978
rect 363498 21922 363554 21978
rect 363622 21922 363678 21978
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 366970 514294 367026 514350
rect 367094 514294 367150 514350
rect 367218 514294 367274 514350
rect 367342 514294 367398 514350
rect 366970 514170 367026 514226
rect 367094 514170 367150 514226
rect 367218 514170 367274 514226
rect 367342 514170 367398 514226
rect 366970 514046 367026 514102
rect 367094 514046 367150 514102
rect 367218 514046 367274 514102
rect 367342 514046 367398 514102
rect 366970 513922 367026 513978
rect 367094 513922 367150 513978
rect 367218 513922 367274 513978
rect 367342 513922 367398 513978
rect 366970 496294 367026 496350
rect 367094 496294 367150 496350
rect 367218 496294 367274 496350
rect 367342 496294 367398 496350
rect 366970 496170 367026 496226
rect 367094 496170 367150 496226
rect 367218 496170 367274 496226
rect 367342 496170 367398 496226
rect 366970 496046 367026 496102
rect 367094 496046 367150 496102
rect 367218 496046 367274 496102
rect 367342 496046 367398 496102
rect 366970 495922 367026 495978
rect 367094 495922 367150 495978
rect 367218 495922 367274 495978
rect 367342 495922 367398 495978
rect 366970 478294 367026 478350
rect 367094 478294 367150 478350
rect 367218 478294 367274 478350
rect 367342 478294 367398 478350
rect 366970 478170 367026 478226
rect 367094 478170 367150 478226
rect 367218 478170 367274 478226
rect 367342 478170 367398 478226
rect 366970 478046 367026 478102
rect 367094 478046 367150 478102
rect 367218 478046 367274 478102
rect 367342 478046 367398 478102
rect 366970 477922 367026 477978
rect 367094 477922 367150 477978
rect 367218 477922 367274 477978
rect 367342 477922 367398 477978
rect 366970 460294 367026 460350
rect 367094 460294 367150 460350
rect 367218 460294 367274 460350
rect 367342 460294 367398 460350
rect 366970 460170 367026 460226
rect 367094 460170 367150 460226
rect 367218 460170 367274 460226
rect 367342 460170 367398 460226
rect 366970 460046 367026 460102
rect 367094 460046 367150 460102
rect 367218 460046 367274 460102
rect 367342 460046 367398 460102
rect 366970 459922 367026 459978
rect 367094 459922 367150 459978
rect 367218 459922 367274 459978
rect 367342 459922 367398 459978
rect 366970 442294 367026 442350
rect 367094 442294 367150 442350
rect 367218 442294 367274 442350
rect 367342 442294 367398 442350
rect 366970 442170 367026 442226
rect 367094 442170 367150 442226
rect 367218 442170 367274 442226
rect 367342 442170 367398 442226
rect 366970 442046 367026 442102
rect 367094 442046 367150 442102
rect 367218 442046 367274 442102
rect 367342 442046 367398 442102
rect 366970 441922 367026 441978
rect 367094 441922 367150 441978
rect 367218 441922 367274 441978
rect 367342 441922 367398 441978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 381250 526294 381306 526350
rect 381374 526294 381430 526350
rect 381498 526294 381554 526350
rect 381622 526294 381678 526350
rect 381250 526170 381306 526226
rect 381374 526170 381430 526226
rect 381498 526170 381554 526226
rect 381622 526170 381678 526226
rect 381250 526046 381306 526102
rect 381374 526046 381430 526102
rect 381498 526046 381554 526102
rect 381622 526046 381678 526102
rect 381250 525922 381306 525978
rect 381374 525922 381430 525978
rect 381498 525922 381554 525978
rect 381622 525922 381678 525978
rect 381250 508294 381306 508350
rect 381374 508294 381430 508350
rect 381498 508294 381554 508350
rect 381622 508294 381678 508350
rect 381250 508170 381306 508226
rect 381374 508170 381430 508226
rect 381498 508170 381554 508226
rect 381622 508170 381678 508226
rect 381250 508046 381306 508102
rect 381374 508046 381430 508102
rect 381498 508046 381554 508102
rect 381622 508046 381678 508102
rect 381250 507922 381306 507978
rect 381374 507922 381430 507978
rect 381498 507922 381554 507978
rect 381622 507922 381678 507978
rect 381250 490294 381306 490350
rect 381374 490294 381430 490350
rect 381498 490294 381554 490350
rect 381622 490294 381678 490350
rect 381250 490170 381306 490226
rect 381374 490170 381430 490226
rect 381498 490170 381554 490226
rect 381622 490170 381678 490226
rect 381250 490046 381306 490102
rect 381374 490046 381430 490102
rect 381498 490046 381554 490102
rect 381622 490046 381678 490102
rect 381250 489922 381306 489978
rect 381374 489922 381430 489978
rect 381498 489922 381554 489978
rect 381622 489922 381678 489978
rect 381250 472294 381306 472350
rect 381374 472294 381430 472350
rect 381498 472294 381554 472350
rect 381622 472294 381678 472350
rect 381250 472170 381306 472226
rect 381374 472170 381430 472226
rect 381498 472170 381554 472226
rect 381622 472170 381678 472226
rect 381250 472046 381306 472102
rect 381374 472046 381430 472102
rect 381498 472046 381554 472102
rect 381622 472046 381678 472102
rect 381250 471922 381306 471978
rect 381374 471922 381430 471978
rect 381498 471922 381554 471978
rect 381622 471922 381678 471978
rect 381250 454294 381306 454350
rect 381374 454294 381430 454350
rect 381498 454294 381554 454350
rect 381622 454294 381678 454350
rect 381250 454170 381306 454226
rect 381374 454170 381430 454226
rect 381498 454170 381554 454226
rect 381622 454170 381678 454226
rect 381250 454046 381306 454102
rect 381374 454046 381430 454102
rect 381498 454046 381554 454102
rect 381622 454046 381678 454102
rect 381250 453922 381306 453978
rect 381374 453922 381430 453978
rect 381498 453922 381554 453978
rect 381622 453922 381678 453978
rect 371718 436261 371774 436317
rect 371842 436261 371898 436317
rect 371718 436137 371774 436193
rect 371842 436137 371898 436193
rect 371718 436013 371774 436069
rect 371842 436013 371898 436069
rect 371718 435889 371774 435945
rect 371842 435889 371898 435945
rect 381250 436294 381306 436350
rect 381374 436294 381430 436350
rect 381498 436294 381554 436350
rect 381622 436294 381678 436350
rect 381250 436170 381306 436226
rect 381374 436170 381430 436226
rect 381498 436170 381554 436226
rect 381622 436170 381678 436226
rect 381250 436046 381306 436102
rect 381374 436046 381430 436102
rect 381498 436046 381554 436102
rect 381622 436046 381678 436102
rect 381250 435922 381306 435978
rect 381374 435922 381430 435978
rect 381498 435922 381554 435978
rect 381622 435922 381678 435978
rect 366970 424294 367026 424350
rect 367094 424294 367150 424350
rect 367218 424294 367274 424350
rect 367342 424294 367398 424350
rect 366970 424170 367026 424226
rect 367094 424170 367150 424226
rect 367218 424170 367274 424226
rect 367342 424170 367398 424226
rect 366970 424046 367026 424102
rect 367094 424046 367150 424102
rect 367218 424046 367274 424102
rect 367342 424046 367398 424102
rect 366970 423922 367026 423978
rect 367094 423922 367150 423978
rect 367218 423922 367274 423978
rect 367342 423922 367398 423978
rect 371718 418294 371774 418350
rect 371842 418294 371898 418350
rect 371718 418170 371774 418226
rect 371842 418170 371898 418226
rect 371718 418046 371774 418102
rect 371842 418046 371898 418102
rect 371718 417922 371774 417978
rect 371842 417922 371898 417978
rect 381250 418294 381306 418350
rect 381374 418294 381430 418350
rect 381498 418294 381554 418350
rect 381622 418294 381678 418350
rect 381250 418170 381306 418226
rect 381374 418170 381430 418226
rect 381498 418170 381554 418226
rect 381622 418170 381678 418226
rect 381250 418046 381306 418102
rect 381374 418046 381430 418102
rect 381498 418046 381554 418102
rect 381622 418046 381678 418102
rect 381250 417922 381306 417978
rect 381374 417922 381430 417978
rect 381498 417922 381554 417978
rect 381622 417922 381678 417978
rect 366970 406294 367026 406350
rect 367094 406294 367150 406350
rect 367218 406294 367274 406350
rect 367342 406294 367398 406350
rect 366970 406170 367026 406226
rect 367094 406170 367150 406226
rect 367218 406170 367274 406226
rect 367342 406170 367398 406226
rect 366970 406046 367026 406102
rect 367094 406046 367150 406102
rect 367218 406046 367274 406102
rect 367342 406046 367398 406102
rect 366970 405922 367026 405978
rect 367094 405922 367150 405978
rect 367218 405922 367274 405978
rect 367342 405922 367398 405978
rect 371718 400294 371774 400350
rect 371842 400294 371898 400350
rect 371718 400170 371774 400226
rect 371842 400170 371898 400226
rect 371718 400046 371774 400102
rect 371842 400046 371898 400102
rect 371718 399922 371774 399978
rect 371842 399922 371898 399978
rect 381250 400294 381306 400350
rect 381374 400294 381430 400350
rect 381498 400294 381554 400350
rect 381622 400294 381678 400350
rect 381250 400170 381306 400226
rect 381374 400170 381430 400226
rect 381498 400170 381554 400226
rect 381622 400170 381678 400226
rect 381250 400046 381306 400102
rect 381374 400046 381430 400102
rect 381498 400046 381554 400102
rect 381622 400046 381678 400102
rect 381250 399922 381306 399978
rect 381374 399922 381430 399978
rect 381498 399922 381554 399978
rect 381622 399922 381678 399978
rect 366970 388294 367026 388350
rect 367094 388294 367150 388350
rect 367218 388294 367274 388350
rect 367342 388294 367398 388350
rect 366970 388170 367026 388226
rect 367094 388170 367150 388226
rect 367218 388170 367274 388226
rect 367342 388170 367398 388226
rect 366970 388046 367026 388102
rect 367094 388046 367150 388102
rect 367218 388046 367274 388102
rect 367342 388046 367398 388102
rect 366970 387922 367026 387978
rect 367094 387922 367150 387978
rect 367218 387922 367274 387978
rect 367342 387922 367398 387978
rect 371718 382294 371774 382350
rect 371842 382294 371898 382350
rect 371718 382170 371774 382226
rect 371842 382170 371898 382226
rect 371718 382046 371774 382102
rect 371842 382046 371898 382102
rect 371718 381922 371774 381978
rect 371842 381922 371898 381978
rect 381250 382294 381306 382350
rect 381374 382294 381430 382350
rect 381498 382294 381554 382350
rect 381622 382294 381678 382350
rect 381250 382170 381306 382226
rect 381374 382170 381430 382226
rect 381498 382170 381554 382226
rect 381622 382170 381678 382226
rect 381250 382046 381306 382102
rect 381374 382046 381430 382102
rect 381498 382046 381554 382102
rect 381622 382046 381678 382102
rect 381250 381922 381306 381978
rect 381374 381922 381430 381978
rect 381498 381922 381554 381978
rect 381622 381922 381678 381978
rect 366970 370294 367026 370350
rect 367094 370294 367150 370350
rect 367218 370294 367274 370350
rect 367342 370294 367398 370350
rect 366970 370170 367026 370226
rect 367094 370170 367150 370226
rect 367218 370170 367274 370226
rect 367342 370170 367398 370226
rect 366970 370046 367026 370102
rect 367094 370046 367150 370102
rect 367218 370046 367274 370102
rect 367342 370046 367398 370102
rect 366970 369922 367026 369978
rect 367094 369922 367150 369978
rect 367218 369922 367274 369978
rect 367342 369922 367398 369978
rect 371718 364294 371774 364350
rect 371842 364294 371898 364350
rect 371718 364170 371774 364226
rect 371842 364170 371898 364226
rect 371718 364046 371774 364102
rect 371842 364046 371898 364102
rect 371718 363922 371774 363978
rect 371842 363922 371898 363978
rect 381250 364294 381306 364350
rect 381374 364294 381430 364350
rect 381498 364294 381554 364350
rect 381622 364294 381678 364350
rect 381250 364170 381306 364226
rect 381374 364170 381430 364226
rect 381498 364170 381554 364226
rect 381622 364170 381678 364226
rect 381250 364046 381306 364102
rect 381374 364046 381430 364102
rect 381498 364046 381554 364102
rect 381622 364046 381678 364102
rect 381250 363922 381306 363978
rect 381374 363922 381430 363978
rect 381498 363922 381554 363978
rect 381622 363922 381678 363978
rect 366970 352294 367026 352350
rect 367094 352294 367150 352350
rect 367218 352294 367274 352350
rect 367342 352294 367398 352350
rect 366970 352170 367026 352226
rect 367094 352170 367150 352226
rect 367218 352170 367274 352226
rect 367342 352170 367398 352226
rect 366970 352046 367026 352102
rect 367094 352046 367150 352102
rect 367218 352046 367274 352102
rect 367342 352046 367398 352102
rect 366970 351922 367026 351978
rect 367094 351922 367150 351978
rect 367218 351922 367274 351978
rect 367342 351922 367398 351978
rect 371718 346294 371774 346350
rect 371842 346294 371898 346350
rect 371718 346170 371774 346226
rect 371842 346170 371898 346226
rect 371718 346046 371774 346102
rect 371842 346046 371898 346102
rect 371718 345922 371774 345978
rect 371842 345922 371898 345978
rect 381250 346294 381306 346350
rect 381374 346294 381430 346350
rect 381498 346294 381554 346350
rect 381622 346294 381678 346350
rect 381250 346170 381306 346226
rect 381374 346170 381430 346226
rect 381498 346170 381554 346226
rect 381622 346170 381678 346226
rect 381250 346046 381306 346102
rect 381374 346046 381430 346102
rect 381498 346046 381554 346102
rect 381622 346046 381678 346102
rect 381250 345922 381306 345978
rect 381374 345922 381430 345978
rect 381498 345922 381554 345978
rect 381622 345922 381678 345978
rect 366970 334294 367026 334350
rect 367094 334294 367150 334350
rect 367218 334294 367274 334350
rect 367342 334294 367398 334350
rect 366970 334170 367026 334226
rect 367094 334170 367150 334226
rect 367218 334170 367274 334226
rect 367342 334170 367398 334226
rect 366970 334046 367026 334102
rect 367094 334046 367150 334102
rect 367218 334046 367274 334102
rect 367342 334046 367398 334102
rect 366970 333922 367026 333978
rect 367094 333922 367150 333978
rect 367218 333922 367274 333978
rect 367342 333922 367398 333978
rect 371718 328294 371774 328350
rect 371842 328294 371898 328350
rect 371718 328170 371774 328226
rect 371842 328170 371898 328226
rect 371718 328046 371774 328102
rect 371842 328046 371898 328102
rect 371718 327922 371774 327978
rect 371842 327922 371898 327978
rect 381250 328294 381306 328350
rect 381374 328294 381430 328350
rect 381498 328294 381554 328350
rect 381622 328294 381678 328350
rect 381250 328170 381306 328226
rect 381374 328170 381430 328226
rect 381498 328170 381554 328226
rect 381622 328170 381678 328226
rect 381250 328046 381306 328102
rect 381374 328046 381430 328102
rect 381498 328046 381554 328102
rect 381622 328046 381678 328102
rect 381250 327922 381306 327978
rect 381374 327922 381430 327978
rect 381498 327922 381554 327978
rect 381622 327922 381678 327978
rect 366970 316294 367026 316350
rect 367094 316294 367150 316350
rect 367218 316294 367274 316350
rect 367342 316294 367398 316350
rect 366970 316170 367026 316226
rect 367094 316170 367150 316226
rect 367218 316170 367274 316226
rect 367342 316170 367398 316226
rect 366970 316046 367026 316102
rect 367094 316046 367150 316102
rect 367218 316046 367274 316102
rect 367342 316046 367398 316102
rect 366970 315922 367026 315978
rect 367094 315922 367150 315978
rect 367218 315922 367274 315978
rect 367342 315922 367398 315978
rect 371718 310294 371774 310350
rect 371842 310294 371898 310350
rect 371718 310170 371774 310226
rect 371842 310170 371898 310226
rect 371718 310046 371774 310102
rect 371842 310046 371898 310102
rect 371718 309922 371774 309978
rect 371842 309922 371898 309978
rect 381250 310294 381306 310350
rect 381374 310294 381430 310350
rect 381498 310294 381554 310350
rect 381622 310294 381678 310350
rect 381250 310170 381306 310226
rect 381374 310170 381430 310226
rect 381498 310170 381554 310226
rect 381622 310170 381678 310226
rect 381250 310046 381306 310102
rect 381374 310046 381430 310102
rect 381498 310046 381554 310102
rect 381622 310046 381678 310102
rect 381250 309922 381306 309978
rect 381374 309922 381430 309978
rect 381498 309922 381554 309978
rect 381622 309922 381678 309978
rect 366970 298294 367026 298350
rect 367094 298294 367150 298350
rect 367218 298294 367274 298350
rect 367342 298294 367398 298350
rect 366970 298170 367026 298226
rect 367094 298170 367150 298226
rect 367218 298170 367274 298226
rect 367342 298170 367398 298226
rect 366970 298046 367026 298102
rect 367094 298046 367150 298102
rect 367218 298046 367274 298102
rect 367342 298046 367398 298102
rect 366970 297922 367026 297978
rect 367094 297922 367150 297978
rect 367218 297922 367274 297978
rect 367342 297922 367398 297978
rect 371718 292294 371774 292350
rect 371842 292294 371898 292350
rect 371718 292170 371774 292226
rect 371842 292170 371898 292226
rect 371718 292046 371774 292102
rect 371842 292046 371898 292102
rect 371718 291922 371774 291978
rect 371842 291922 371898 291978
rect 381250 292294 381306 292350
rect 381374 292294 381430 292350
rect 381498 292294 381554 292350
rect 381622 292294 381678 292350
rect 381250 292170 381306 292226
rect 381374 292170 381430 292226
rect 381498 292170 381554 292226
rect 381622 292170 381678 292226
rect 381250 292046 381306 292102
rect 381374 292046 381430 292102
rect 381498 292046 381554 292102
rect 381622 292046 381678 292102
rect 381250 291922 381306 291978
rect 381374 291922 381430 291978
rect 381498 291922 381554 291978
rect 381622 291922 381678 291978
rect 366970 280294 367026 280350
rect 367094 280294 367150 280350
rect 367218 280294 367274 280350
rect 367342 280294 367398 280350
rect 366970 280170 367026 280226
rect 367094 280170 367150 280226
rect 367218 280170 367274 280226
rect 367342 280170 367398 280226
rect 366970 280046 367026 280102
rect 367094 280046 367150 280102
rect 367218 280046 367274 280102
rect 367342 280046 367398 280102
rect 366970 279922 367026 279978
rect 367094 279922 367150 279978
rect 367218 279922 367274 279978
rect 367342 279922 367398 279978
rect 371718 274294 371774 274350
rect 371842 274294 371898 274350
rect 371718 274170 371774 274226
rect 371842 274170 371898 274226
rect 371718 274046 371774 274102
rect 371842 274046 371898 274102
rect 371718 273922 371774 273978
rect 371842 273922 371898 273978
rect 381250 274294 381306 274350
rect 381374 274294 381430 274350
rect 381498 274294 381554 274350
rect 381622 274294 381678 274350
rect 381250 274170 381306 274226
rect 381374 274170 381430 274226
rect 381498 274170 381554 274226
rect 381622 274170 381678 274226
rect 381250 274046 381306 274102
rect 381374 274046 381430 274102
rect 381498 274046 381554 274102
rect 381622 274046 381678 274102
rect 381250 273922 381306 273978
rect 381374 273922 381430 273978
rect 381498 273922 381554 273978
rect 381622 273922 381678 273978
rect 366970 262294 367026 262350
rect 367094 262294 367150 262350
rect 367218 262294 367274 262350
rect 367342 262294 367398 262350
rect 366970 262170 367026 262226
rect 367094 262170 367150 262226
rect 367218 262170 367274 262226
rect 367342 262170 367398 262226
rect 366970 262046 367026 262102
rect 367094 262046 367150 262102
rect 367218 262046 367274 262102
rect 367342 262046 367398 262102
rect 366970 261922 367026 261978
rect 367094 261922 367150 261978
rect 367218 261922 367274 261978
rect 367342 261922 367398 261978
rect 371718 256294 371774 256350
rect 371842 256294 371898 256350
rect 371718 256170 371774 256226
rect 371842 256170 371898 256226
rect 371718 256046 371774 256102
rect 371842 256046 371898 256102
rect 371718 255922 371774 255978
rect 371842 255922 371898 255978
rect 381250 256294 381306 256350
rect 381374 256294 381430 256350
rect 381498 256294 381554 256350
rect 381622 256294 381678 256350
rect 381250 256170 381306 256226
rect 381374 256170 381430 256226
rect 381498 256170 381554 256226
rect 381622 256170 381678 256226
rect 381250 256046 381306 256102
rect 381374 256046 381430 256102
rect 381498 256046 381554 256102
rect 381622 256046 381678 256102
rect 381250 255922 381306 255978
rect 381374 255922 381430 255978
rect 381498 255922 381554 255978
rect 381622 255922 381678 255978
rect 366970 244294 367026 244350
rect 367094 244294 367150 244350
rect 367218 244294 367274 244350
rect 367342 244294 367398 244350
rect 366970 244170 367026 244226
rect 367094 244170 367150 244226
rect 367218 244170 367274 244226
rect 367342 244170 367398 244226
rect 366970 244046 367026 244102
rect 367094 244046 367150 244102
rect 367218 244046 367274 244102
rect 367342 244046 367398 244102
rect 366970 243922 367026 243978
rect 367094 243922 367150 243978
rect 367218 243922 367274 243978
rect 367342 243922 367398 243978
rect 371718 238294 371774 238350
rect 371842 238294 371898 238350
rect 371718 238170 371774 238226
rect 371842 238170 371898 238226
rect 371718 238046 371774 238102
rect 371842 238046 371898 238102
rect 371718 237922 371774 237978
rect 371842 237922 371898 237978
rect 381250 238294 381306 238350
rect 381374 238294 381430 238350
rect 381498 238294 381554 238350
rect 381622 238294 381678 238350
rect 381250 238170 381306 238226
rect 381374 238170 381430 238226
rect 381498 238170 381554 238226
rect 381622 238170 381678 238226
rect 381250 238046 381306 238102
rect 381374 238046 381430 238102
rect 381498 238046 381554 238102
rect 381622 238046 381678 238102
rect 381250 237922 381306 237978
rect 381374 237922 381430 237978
rect 381498 237922 381554 237978
rect 381622 237922 381678 237978
rect 366970 226294 367026 226350
rect 367094 226294 367150 226350
rect 367218 226294 367274 226350
rect 367342 226294 367398 226350
rect 366970 226170 367026 226226
rect 367094 226170 367150 226226
rect 367218 226170 367274 226226
rect 367342 226170 367398 226226
rect 366970 226046 367026 226102
rect 367094 226046 367150 226102
rect 367218 226046 367274 226102
rect 367342 226046 367398 226102
rect 366970 225922 367026 225978
rect 367094 225922 367150 225978
rect 367218 225922 367274 225978
rect 367342 225922 367398 225978
rect 371718 220294 371774 220350
rect 371842 220294 371898 220350
rect 371718 220170 371774 220226
rect 371842 220170 371898 220226
rect 371718 220046 371774 220102
rect 371842 220046 371898 220102
rect 371718 219922 371774 219978
rect 371842 219922 371898 219978
rect 381250 220294 381306 220350
rect 381374 220294 381430 220350
rect 381498 220294 381554 220350
rect 381622 220294 381678 220350
rect 381250 220170 381306 220226
rect 381374 220170 381430 220226
rect 381498 220170 381554 220226
rect 381622 220170 381678 220226
rect 381250 220046 381306 220102
rect 381374 220046 381430 220102
rect 381498 220046 381554 220102
rect 381622 220046 381678 220102
rect 381250 219922 381306 219978
rect 381374 219922 381430 219978
rect 381498 219922 381554 219978
rect 381622 219922 381678 219978
rect 366970 208294 367026 208350
rect 367094 208294 367150 208350
rect 367218 208294 367274 208350
rect 367342 208294 367398 208350
rect 366970 208170 367026 208226
rect 367094 208170 367150 208226
rect 367218 208170 367274 208226
rect 367342 208170 367398 208226
rect 366970 208046 367026 208102
rect 367094 208046 367150 208102
rect 367218 208046 367274 208102
rect 367342 208046 367398 208102
rect 366970 207922 367026 207978
rect 367094 207922 367150 207978
rect 367218 207922 367274 207978
rect 367342 207922 367398 207978
rect 371718 202294 371774 202350
rect 371842 202294 371898 202350
rect 371718 202170 371774 202226
rect 371842 202170 371898 202226
rect 371718 202046 371774 202102
rect 371842 202046 371898 202102
rect 371718 201922 371774 201978
rect 371842 201922 371898 201978
rect 381250 202294 381306 202350
rect 381374 202294 381430 202350
rect 381498 202294 381554 202350
rect 381622 202294 381678 202350
rect 381250 202170 381306 202226
rect 381374 202170 381430 202226
rect 381498 202170 381554 202226
rect 381622 202170 381678 202226
rect 381250 202046 381306 202102
rect 381374 202046 381430 202102
rect 381498 202046 381554 202102
rect 381622 202046 381678 202102
rect 381250 201922 381306 201978
rect 381374 201922 381430 201978
rect 381498 201922 381554 201978
rect 381622 201922 381678 201978
rect 366970 190294 367026 190350
rect 367094 190294 367150 190350
rect 367218 190294 367274 190350
rect 367342 190294 367398 190350
rect 366970 190170 367026 190226
rect 367094 190170 367150 190226
rect 367218 190170 367274 190226
rect 367342 190170 367398 190226
rect 366970 190046 367026 190102
rect 367094 190046 367150 190102
rect 367218 190046 367274 190102
rect 367342 190046 367398 190102
rect 366970 189922 367026 189978
rect 367094 189922 367150 189978
rect 367218 189922 367274 189978
rect 367342 189922 367398 189978
rect 371718 184294 371774 184350
rect 371842 184294 371898 184350
rect 371718 184170 371774 184226
rect 371842 184170 371898 184226
rect 371718 184046 371774 184102
rect 371842 184046 371898 184102
rect 371718 183922 371774 183978
rect 371842 183922 371898 183978
rect 381250 184294 381306 184350
rect 381374 184294 381430 184350
rect 381498 184294 381554 184350
rect 381622 184294 381678 184350
rect 381250 184170 381306 184226
rect 381374 184170 381430 184226
rect 381498 184170 381554 184226
rect 381622 184170 381678 184226
rect 381250 184046 381306 184102
rect 381374 184046 381430 184102
rect 381498 184046 381554 184102
rect 381622 184046 381678 184102
rect 381250 183922 381306 183978
rect 381374 183922 381430 183978
rect 381498 183922 381554 183978
rect 381622 183922 381678 183978
rect 366970 172294 367026 172350
rect 367094 172294 367150 172350
rect 367218 172294 367274 172350
rect 367342 172294 367398 172350
rect 366970 172170 367026 172226
rect 367094 172170 367150 172226
rect 367218 172170 367274 172226
rect 367342 172170 367398 172226
rect 366970 172046 367026 172102
rect 367094 172046 367150 172102
rect 367218 172046 367274 172102
rect 367342 172046 367398 172102
rect 366970 171922 367026 171978
rect 367094 171922 367150 171978
rect 367218 171922 367274 171978
rect 367342 171922 367398 171978
rect 371718 166294 371774 166350
rect 371842 166294 371898 166350
rect 371718 166170 371774 166226
rect 371842 166170 371898 166226
rect 371718 166046 371774 166102
rect 371842 166046 371898 166102
rect 371718 165922 371774 165978
rect 371842 165922 371898 165978
rect 381250 166294 381306 166350
rect 381374 166294 381430 166350
rect 381498 166294 381554 166350
rect 381622 166294 381678 166350
rect 381250 166170 381306 166226
rect 381374 166170 381430 166226
rect 381498 166170 381554 166226
rect 381622 166170 381678 166226
rect 381250 166046 381306 166102
rect 381374 166046 381430 166102
rect 381498 166046 381554 166102
rect 381622 166046 381678 166102
rect 381250 165922 381306 165978
rect 381374 165922 381430 165978
rect 381498 165922 381554 165978
rect 381622 165922 381678 165978
rect 366970 154294 367026 154350
rect 367094 154294 367150 154350
rect 367218 154294 367274 154350
rect 367342 154294 367398 154350
rect 366970 154170 367026 154226
rect 367094 154170 367150 154226
rect 367218 154170 367274 154226
rect 367342 154170 367398 154226
rect 366970 154046 367026 154102
rect 367094 154046 367150 154102
rect 367218 154046 367274 154102
rect 367342 154046 367398 154102
rect 366970 153922 367026 153978
rect 367094 153922 367150 153978
rect 367218 153922 367274 153978
rect 367342 153922 367398 153978
rect 371718 148294 371774 148350
rect 371842 148294 371898 148350
rect 371718 148170 371774 148226
rect 371842 148170 371898 148226
rect 371718 148046 371774 148102
rect 371842 148046 371898 148102
rect 371718 147922 371774 147978
rect 371842 147922 371898 147978
rect 381250 148294 381306 148350
rect 381374 148294 381430 148350
rect 381498 148294 381554 148350
rect 381622 148294 381678 148350
rect 381250 148170 381306 148226
rect 381374 148170 381430 148226
rect 381498 148170 381554 148226
rect 381622 148170 381678 148226
rect 381250 148046 381306 148102
rect 381374 148046 381430 148102
rect 381498 148046 381554 148102
rect 381622 148046 381678 148102
rect 381250 147922 381306 147978
rect 381374 147922 381430 147978
rect 381498 147922 381554 147978
rect 381622 147922 381678 147978
rect 366970 136294 367026 136350
rect 367094 136294 367150 136350
rect 367218 136294 367274 136350
rect 367342 136294 367398 136350
rect 366970 136170 367026 136226
rect 367094 136170 367150 136226
rect 367218 136170 367274 136226
rect 367342 136170 367398 136226
rect 366970 136046 367026 136102
rect 367094 136046 367150 136102
rect 367218 136046 367274 136102
rect 367342 136046 367398 136102
rect 366970 135922 367026 135978
rect 367094 135922 367150 135978
rect 367218 135922 367274 135978
rect 367342 135922 367398 135978
rect 371718 130294 371774 130350
rect 371842 130294 371898 130350
rect 371718 130170 371774 130226
rect 371842 130170 371898 130226
rect 371718 130046 371774 130102
rect 371842 130046 371898 130102
rect 371718 129922 371774 129978
rect 371842 129922 371898 129978
rect 381250 130294 381306 130350
rect 381374 130294 381430 130350
rect 381498 130294 381554 130350
rect 381622 130294 381678 130350
rect 381250 130170 381306 130226
rect 381374 130170 381430 130226
rect 381498 130170 381554 130226
rect 381622 130170 381678 130226
rect 381250 130046 381306 130102
rect 381374 130046 381430 130102
rect 381498 130046 381554 130102
rect 381622 130046 381678 130102
rect 381250 129922 381306 129978
rect 381374 129922 381430 129978
rect 381498 129922 381554 129978
rect 381622 129922 381678 129978
rect 366970 118294 367026 118350
rect 367094 118294 367150 118350
rect 367218 118294 367274 118350
rect 367342 118294 367398 118350
rect 366970 118170 367026 118226
rect 367094 118170 367150 118226
rect 367218 118170 367274 118226
rect 367342 118170 367398 118226
rect 366970 118046 367026 118102
rect 367094 118046 367150 118102
rect 367218 118046 367274 118102
rect 367342 118046 367398 118102
rect 366970 117922 367026 117978
rect 367094 117922 367150 117978
rect 367218 117922 367274 117978
rect 367342 117922 367398 117978
rect 371718 112294 371774 112350
rect 371842 112294 371898 112350
rect 371718 112170 371774 112226
rect 371842 112170 371898 112226
rect 371718 112046 371774 112102
rect 371842 112046 371898 112102
rect 371718 111922 371774 111978
rect 371842 111922 371898 111978
rect 381250 112294 381306 112350
rect 381374 112294 381430 112350
rect 381498 112294 381554 112350
rect 381622 112294 381678 112350
rect 381250 112170 381306 112226
rect 381374 112170 381430 112226
rect 381498 112170 381554 112226
rect 381622 112170 381678 112226
rect 381250 112046 381306 112102
rect 381374 112046 381430 112102
rect 381498 112046 381554 112102
rect 381622 112046 381678 112102
rect 381250 111922 381306 111978
rect 381374 111922 381430 111978
rect 381498 111922 381554 111978
rect 381622 111922 381678 111978
rect 366970 100294 367026 100350
rect 367094 100294 367150 100350
rect 367218 100294 367274 100350
rect 367342 100294 367398 100350
rect 366970 100170 367026 100226
rect 367094 100170 367150 100226
rect 367218 100170 367274 100226
rect 367342 100170 367398 100226
rect 366970 100046 367026 100102
rect 367094 100046 367150 100102
rect 367218 100046 367274 100102
rect 367342 100046 367398 100102
rect 366970 99922 367026 99978
rect 367094 99922 367150 99978
rect 367218 99922 367274 99978
rect 367342 99922 367398 99978
rect 371718 94294 371774 94350
rect 371842 94294 371898 94350
rect 371718 94170 371774 94226
rect 371842 94170 371898 94226
rect 371718 94046 371774 94102
rect 371842 94046 371898 94102
rect 371718 93922 371774 93978
rect 371842 93922 371898 93978
rect 381250 94294 381306 94350
rect 381374 94294 381430 94350
rect 381498 94294 381554 94350
rect 381622 94294 381678 94350
rect 381250 94170 381306 94226
rect 381374 94170 381430 94226
rect 381498 94170 381554 94226
rect 381622 94170 381678 94226
rect 381250 94046 381306 94102
rect 381374 94046 381430 94102
rect 381498 94046 381554 94102
rect 381622 94046 381678 94102
rect 381250 93922 381306 93978
rect 381374 93922 381430 93978
rect 381498 93922 381554 93978
rect 381622 93922 381678 93978
rect 366970 82294 367026 82350
rect 367094 82294 367150 82350
rect 367218 82294 367274 82350
rect 367342 82294 367398 82350
rect 366970 82170 367026 82226
rect 367094 82170 367150 82226
rect 367218 82170 367274 82226
rect 367342 82170 367398 82226
rect 366970 82046 367026 82102
rect 367094 82046 367150 82102
rect 367218 82046 367274 82102
rect 367342 82046 367398 82102
rect 366970 81922 367026 81978
rect 367094 81922 367150 81978
rect 367218 81922 367274 81978
rect 367342 81922 367398 81978
rect 371718 76294 371774 76350
rect 371842 76294 371898 76350
rect 371718 76170 371774 76226
rect 371842 76170 371898 76226
rect 371718 76046 371774 76102
rect 371842 76046 371898 76102
rect 371718 75922 371774 75978
rect 371842 75922 371898 75978
rect 381250 76294 381306 76350
rect 381374 76294 381430 76350
rect 381498 76294 381554 76350
rect 381622 76294 381678 76350
rect 381250 76170 381306 76226
rect 381374 76170 381430 76226
rect 381498 76170 381554 76226
rect 381622 76170 381678 76226
rect 381250 76046 381306 76102
rect 381374 76046 381430 76102
rect 381498 76046 381554 76102
rect 381622 76046 381678 76102
rect 381250 75922 381306 75978
rect 381374 75922 381430 75978
rect 381498 75922 381554 75978
rect 381622 75922 381678 75978
rect 366970 64294 367026 64350
rect 367094 64294 367150 64350
rect 367218 64294 367274 64350
rect 367342 64294 367398 64350
rect 366970 64170 367026 64226
rect 367094 64170 367150 64226
rect 367218 64170 367274 64226
rect 367342 64170 367398 64226
rect 366970 64046 367026 64102
rect 367094 64046 367150 64102
rect 367218 64046 367274 64102
rect 367342 64046 367398 64102
rect 366970 63922 367026 63978
rect 367094 63922 367150 63978
rect 367218 63922 367274 63978
rect 367342 63922 367398 63978
rect 366970 46294 367026 46350
rect 367094 46294 367150 46350
rect 367218 46294 367274 46350
rect 367342 46294 367398 46350
rect 366970 46170 367026 46226
rect 367094 46170 367150 46226
rect 367218 46170 367274 46226
rect 367342 46170 367398 46226
rect 366970 46046 367026 46102
rect 367094 46046 367150 46102
rect 367218 46046 367274 46102
rect 367342 46046 367398 46102
rect 366970 45922 367026 45978
rect 367094 45922 367150 45978
rect 367218 45922 367274 45978
rect 367342 45922 367398 45978
rect 366970 28294 367026 28350
rect 367094 28294 367150 28350
rect 367218 28294 367274 28350
rect 367342 28294 367398 28350
rect 366970 28170 367026 28226
rect 367094 28170 367150 28226
rect 367218 28170 367274 28226
rect 367342 28170 367398 28226
rect 366970 28046 367026 28102
rect 367094 28046 367150 28102
rect 367218 28046 367274 28102
rect 367342 28046 367398 28102
rect 366970 27922 367026 27978
rect 367094 27922 367150 27978
rect 367218 27922 367274 27978
rect 367342 27922 367398 27978
rect 366970 10294 367026 10350
rect 367094 10294 367150 10350
rect 367218 10294 367274 10350
rect 367342 10294 367398 10350
rect 366970 10170 367026 10226
rect 367094 10170 367150 10226
rect 367218 10170 367274 10226
rect 367342 10170 367398 10226
rect 366970 10046 367026 10102
rect 367094 10046 367150 10102
rect 367218 10046 367274 10102
rect 367342 10046 367398 10102
rect 366970 9922 367026 9978
rect 367094 9922 367150 9978
rect 367218 9922 367274 9978
rect 367342 9922 367398 9978
rect 366970 -1176 367026 -1120
rect 367094 -1176 367150 -1120
rect 367218 -1176 367274 -1120
rect 367342 -1176 367398 -1120
rect 366970 -1300 367026 -1244
rect 367094 -1300 367150 -1244
rect 367218 -1300 367274 -1244
rect 367342 -1300 367398 -1244
rect 366970 -1424 367026 -1368
rect 367094 -1424 367150 -1368
rect 367218 -1424 367274 -1368
rect 367342 -1424 367398 -1368
rect 366970 -1548 367026 -1492
rect 367094 -1548 367150 -1492
rect 367218 -1548 367274 -1492
rect 367342 -1548 367398 -1492
rect 381250 58294 381306 58350
rect 381374 58294 381430 58350
rect 381498 58294 381554 58350
rect 381622 58294 381678 58350
rect 381250 58170 381306 58226
rect 381374 58170 381430 58226
rect 381498 58170 381554 58226
rect 381622 58170 381678 58226
rect 381250 58046 381306 58102
rect 381374 58046 381430 58102
rect 381498 58046 381554 58102
rect 381622 58046 381678 58102
rect 381250 57922 381306 57978
rect 381374 57922 381430 57978
rect 381498 57922 381554 57978
rect 381622 57922 381678 57978
rect 381250 40294 381306 40350
rect 381374 40294 381430 40350
rect 381498 40294 381554 40350
rect 381622 40294 381678 40350
rect 381250 40170 381306 40226
rect 381374 40170 381430 40226
rect 381498 40170 381554 40226
rect 381622 40170 381678 40226
rect 381250 40046 381306 40102
rect 381374 40046 381430 40102
rect 381498 40046 381554 40102
rect 381622 40046 381678 40102
rect 381250 39922 381306 39978
rect 381374 39922 381430 39978
rect 381498 39922 381554 39978
rect 381622 39922 381678 39978
rect 381250 22294 381306 22350
rect 381374 22294 381430 22350
rect 381498 22294 381554 22350
rect 381622 22294 381678 22350
rect 381250 22170 381306 22226
rect 381374 22170 381430 22226
rect 381498 22170 381554 22226
rect 381622 22170 381678 22226
rect 381250 22046 381306 22102
rect 381374 22046 381430 22102
rect 381498 22046 381554 22102
rect 381622 22046 381678 22102
rect 381250 21922 381306 21978
rect 381374 21922 381430 21978
rect 381498 21922 381554 21978
rect 381622 21922 381678 21978
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 598116 385026 598172
rect 385094 598116 385150 598172
rect 385218 598116 385274 598172
rect 385342 598116 385398 598172
rect 384970 597992 385026 598048
rect 385094 597992 385150 598048
rect 385218 597992 385274 598048
rect 385342 597992 385398 598048
rect 384970 597868 385026 597924
rect 385094 597868 385150 597924
rect 385218 597868 385274 597924
rect 385342 597868 385398 597924
rect 384970 597744 385026 597800
rect 385094 597744 385150 597800
rect 385218 597744 385274 597800
rect 385342 597744 385398 597800
rect 384970 586294 385026 586350
rect 385094 586294 385150 586350
rect 385218 586294 385274 586350
rect 385342 586294 385398 586350
rect 384970 586170 385026 586226
rect 385094 586170 385150 586226
rect 385218 586170 385274 586226
rect 385342 586170 385398 586226
rect 384970 586046 385026 586102
rect 385094 586046 385150 586102
rect 385218 586046 385274 586102
rect 385342 586046 385398 586102
rect 384970 585922 385026 585978
rect 385094 585922 385150 585978
rect 385218 585922 385274 585978
rect 385342 585922 385398 585978
rect 384970 568294 385026 568350
rect 385094 568294 385150 568350
rect 385218 568294 385274 568350
rect 385342 568294 385398 568350
rect 384970 568170 385026 568226
rect 385094 568170 385150 568226
rect 385218 568170 385274 568226
rect 385342 568170 385398 568226
rect 384970 568046 385026 568102
rect 385094 568046 385150 568102
rect 385218 568046 385274 568102
rect 385342 568046 385398 568102
rect 384970 567922 385026 567978
rect 385094 567922 385150 567978
rect 385218 567922 385274 567978
rect 385342 567922 385398 567978
rect 384970 550294 385026 550350
rect 385094 550294 385150 550350
rect 385218 550294 385274 550350
rect 385342 550294 385398 550350
rect 384970 550170 385026 550226
rect 385094 550170 385150 550226
rect 385218 550170 385274 550226
rect 385342 550170 385398 550226
rect 384970 550046 385026 550102
rect 385094 550046 385150 550102
rect 385218 550046 385274 550102
rect 385342 550046 385398 550102
rect 384970 549922 385026 549978
rect 385094 549922 385150 549978
rect 385218 549922 385274 549978
rect 385342 549922 385398 549978
rect 384970 532294 385026 532350
rect 385094 532294 385150 532350
rect 385218 532294 385274 532350
rect 385342 532294 385398 532350
rect 384970 532170 385026 532226
rect 385094 532170 385150 532226
rect 385218 532170 385274 532226
rect 385342 532170 385398 532226
rect 384970 532046 385026 532102
rect 385094 532046 385150 532102
rect 385218 532046 385274 532102
rect 385342 532046 385398 532102
rect 384970 531922 385026 531978
rect 385094 531922 385150 531978
rect 385218 531922 385274 531978
rect 385342 531922 385398 531978
rect 384970 514294 385026 514350
rect 385094 514294 385150 514350
rect 385218 514294 385274 514350
rect 385342 514294 385398 514350
rect 384970 514170 385026 514226
rect 385094 514170 385150 514226
rect 385218 514170 385274 514226
rect 385342 514170 385398 514226
rect 384970 514046 385026 514102
rect 385094 514046 385150 514102
rect 385218 514046 385274 514102
rect 385342 514046 385398 514102
rect 384970 513922 385026 513978
rect 385094 513922 385150 513978
rect 385218 513922 385274 513978
rect 385342 513922 385398 513978
rect 384970 496294 385026 496350
rect 385094 496294 385150 496350
rect 385218 496294 385274 496350
rect 385342 496294 385398 496350
rect 384970 496170 385026 496226
rect 385094 496170 385150 496226
rect 385218 496170 385274 496226
rect 385342 496170 385398 496226
rect 384970 496046 385026 496102
rect 385094 496046 385150 496102
rect 385218 496046 385274 496102
rect 385342 496046 385398 496102
rect 384970 495922 385026 495978
rect 385094 495922 385150 495978
rect 385218 495922 385274 495978
rect 385342 495922 385398 495978
rect 384970 478294 385026 478350
rect 385094 478294 385150 478350
rect 385218 478294 385274 478350
rect 385342 478294 385398 478350
rect 384970 478170 385026 478226
rect 385094 478170 385150 478226
rect 385218 478170 385274 478226
rect 385342 478170 385398 478226
rect 384970 478046 385026 478102
rect 385094 478046 385150 478102
rect 385218 478046 385274 478102
rect 385342 478046 385398 478102
rect 384970 477922 385026 477978
rect 385094 477922 385150 477978
rect 385218 477922 385274 477978
rect 385342 477922 385398 477978
rect 384970 460294 385026 460350
rect 385094 460294 385150 460350
rect 385218 460294 385274 460350
rect 385342 460294 385398 460350
rect 384970 460170 385026 460226
rect 385094 460170 385150 460226
rect 385218 460170 385274 460226
rect 385342 460170 385398 460226
rect 384970 460046 385026 460102
rect 385094 460046 385150 460102
rect 385218 460046 385274 460102
rect 385342 460046 385398 460102
rect 384970 459922 385026 459978
rect 385094 459922 385150 459978
rect 385218 459922 385274 459978
rect 385342 459922 385398 459978
rect 384970 442294 385026 442350
rect 385094 442294 385150 442350
rect 385218 442294 385274 442350
rect 385342 442294 385398 442350
rect 384970 442170 385026 442226
rect 385094 442170 385150 442226
rect 385218 442170 385274 442226
rect 385342 442170 385398 442226
rect 384970 442046 385026 442102
rect 385094 442046 385150 442102
rect 385218 442046 385274 442102
rect 385342 442046 385398 442102
rect 384970 441922 385026 441978
rect 385094 441922 385150 441978
rect 385218 441922 385274 441978
rect 385342 441922 385398 441978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 399250 526294 399306 526350
rect 399374 526294 399430 526350
rect 399498 526294 399554 526350
rect 399622 526294 399678 526350
rect 399250 526170 399306 526226
rect 399374 526170 399430 526226
rect 399498 526170 399554 526226
rect 399622 526170 399678 526226
rect 399250 526046 399306 526102
rect 399374 526046 399430 526102
rect 399498 526046 399554 526102
rect 399622 526046 399678 526102
rect 399250 525922 399306 525978
rect 399374 525922 399430 525978
rect 399498 525922 399554 525978
rect 399622 525922 399678 525978
rect 399250 508294 399306 508350
rect 399374 508294 399430 508350
rect 399498 508294 399554 508350
rect 399622 508294 399678 508350
rect 399250 508170 399306 508226
rect 399374 508170 399430 508226
rect 399498 508170 399554 508226
rect 399622 508170 399678 508226
rect 399250 508046 399306 508102
rect 399374 508046 399430 508102
rect 399498 508046 399554 508102
rect 399622 508046 399678 508102
rect 399250 507922 399306 507978
rect 399374 507922 399430 507978
rect 399498 507922 399554 507978
rect 399622 507922 399678 507978
rect 399250 490294 399306 490350
rect 399374 490294 399430 490350
rect 399498 490294 399554 490350
rect 399622 490294 399678 490350
rect 399250 490170 399306 490226
rect 399374 490170 399430 490226
rect 399498 490170 399554 490226
rect 399622 490170 399678 490226
rect 399250 490046 399306 490102
rect 399374 490046 399430 490102
rect 399498 490046 399554 490102
rect 399622 490046 399678 490102
rect 399250 489922 399306 489978
rect 399374 489922 399430 489978
rect 399498 489922 399554 489978
rect 399622 489922 399678 489978
rect 399250 472294 399306 472350
rect 399374 472294 399430 472350
rect 399498 472294 399554 472350
rect 399622 472294 399678 472350
rect 399250 472170 399306 472226
rect 399374 472170 399430 472226
rect 399498 472170 399554 472226
rect 399622 472170 399678 472226
rect 399250 472046 399306 472102
rect 399374 472046 399430 472102
rect 399498 472046 399554 472102
rect 399622 472046 399678 472102
rect 399250 471922 399306 471978
rect 399374 471922 399430 471978
rect 399498 471922 399554 471978
rect 399622 471922 399678 471978
rect 399250 454294 399306 454350
rect 399374 454294 399430 454350
rect 399498 454294 399554 454350
rect 399622 454294 399678 454350
rect 399250 454170 399306 454226
rect 399374 454170 399430 454226
rect 399498 454170 399554 454226
rect 399622 454170 399678 454226
rect 399250 454046 399306 454102
rect 399374 454046 399430 454102
rect 399498 454046 399554 454102
rect 399622 454046 399678 454102
rect 399250 453922 399306 453978
rect 399374 453922 399430 453978
rect 399498 453922 399554 453978
rect 399622 453922 399678 453978
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 402970 514294 403026 514350
rect 403094 514294 403150 514350
rect 403218 514294 403274 514350
rect 403342 514294 403398 514350
rect 402970 514170 403026 514226
rect 403094 514170 403150 514226
rect 403218 514170 403274 514226
rect 403342 514170 403398 514226
rect 402970 514046 403026 514102
rect 403094 514046 403150 514102
rect 403218 514046 403274 514102
rect 403342 514046 403398 514102
rect 402970 513922 403026 513978
rect 403094 513922 403150 513978
rect 403218 513922 403274 513978
rect 403342 513922 403398 513978
rect 402970 496294 403026 496350
rect 403094 496294 403150 496350
rect 403218 496294 403274 496350
rect 403342 496294 403398 496350
rect 402970 496170 403026 496226
rect 403094 496170 403150 496226
rect 403218 496170 403274 496226
rect 403342 496170 403398 496226
rect 402970 496046 403026 496102
rect 403094 496046 403150 496102
rect 403218 496046 403274 496102
rect 403342 496046 403398 496102
rect 402970 495922 403026 495978
rect 403094 495922 403150 495978
rect 403218 495922 403274 495978
rect 403342 495922 403398 495978
rect 402970 478294 403026 478350
rect 403094 478294 403150 478350
rect 403218 478294 403274 478350
rect 403342 478294 403398 478350
rect 402970 478170 403026 478226
rect 403094 478170 403150 478226
rect 403218 478170 403274 478226
rect 403342 478170 403398 478226
rect 402970 478046 403026 478102
rect 403094 478046 403150 478102
rect 403218 478046 403274 478102
rect 403342 478046 403398 478102
rect 402970 477922 403026 477978
rect 403094 477922 403150 477978
rect 403218 477922 403274 477978
rect 403342 477922 403398 477978
rect 402970 460294 403026 460350
rect 403094 460294 403150 460350
rect 403218 460294 403274 460350
rect 403342 460294 403398 460350
rect 402970 460170 403026 460226
rect 403094 460170 403150 460226
rect 403218 460170 403274 460226
rect 403342 460170 403398 460226
rect 402970 460046 403026 460102
rect 403094 460046 403150 460102
rect 403218 460046 403274 460102
rect 403342 460046 403398 460102
rect 402970 459922 403026 459978
rect 403094 459922 403150 459978
rect 403218 459922 403274 459978
rect 403342 459922 403398 459978
rect 402970 442294 403026 442350
rect 403094 442294 403150 442350
rect 403218 442294 403274 442350
rect 403342 442294 403398 442350
rect 402970 442170 403026 442226
rect 403094 442170 403150 442226
rect 403218 442170 403274 442226
rect 403342 442170 403398 442226
rect 402970 442046 403026 442102
rect 403094 442046 403150 442102
rect 403218 442046 403274 442102
rect 403342 442046 403398 442102
rect 402970 441922 403026 441978
rect 403094 441922 403150 441978
rect 403218 441922 403274 441978
rect 403342 441922 403398 441978
rect 399250 436294 399306 436350
rect 399374 436294 399430 436350
rect 399498 436294 399554 436350
rect 399622 436294 399678 436350
rect 399250 436170 399306 436226
rect 399374 436170 399430 436226
rect 399498 436170 399554 436226
rect 399622 436170 399678 436226
rect 399250 436046 399306 436102
rect 399374 436046 399430 436102
rect 399498 436046 399554 436102
rect 399622 436046 399678 436102
rect 399250 435922 399306 435978
rect 399374 435922 399430 435978
rect 399498 435922 399554 435978
rect 399622 435922 399678 435978
rect 384970 424294 385026 424350
rect 385094 424294 385150 424350
rect 385218 424294 385274 424350
rect 385342 424294 385398 424350
rect 384970 424170 385026 424226
rect 385094 424170 385150 424226
rect 385218 424170 385274 424226
rect 385342 424170 385398 424226
rect 384970 424046 385026 424102
rect 385094 424046 385150 424102
rect 385218 424046 385274 424102
rect 385342 424046 385398 424102
rect 384970 423922 385026 423978
rect 385094 423922 385150 423978
rect 385218 423922 385274 423978
rect 385342 423922 385398 423978
rect 387078 424294 387134 424350
rect 387202 424294 387258 424350
rect 387078 424170 387134 424226
rect 387202 424170 387258 424226
rect 387078 424046 387134 424102
rect 387202 424046 387258 424102
rect 387078 423922 387134 423978
rect 387202 423922 387258 423978
rect 402438 436261 402494 436317
rect 402562 436261 402618 436317
rect 402438 436137 402494 436193
rect 402562 436137 402618 436193
rect 402438 436013 402494 436069
rect 402562 436013 402618 436069
rect 402438 435889 402494 435945
rect 402562 435889 402618 435945
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 417250 526294 417306 526350
rect 417374 526294 417430 526350
rect 417498 526294 417554 526350
rect 417622 526294 417678 526350
rect 417250 526170 417306 526226
rect 417374 526170 417430 526226
rect 417498 526170 417554 526226
rect 417622 526170 417678 526226
rect 417250 526046 417306 526102
rect 417374 526046 417430 526102
rect 417498 526046 417554 526102
rect 417622 526046 417678 526102
rect 417250 525922 417306 525978
rect 417374 525922 417430 525978
rect 417498 525922 417554 525978
rect 417622 525922 417678 525978
rect 417250 508294 417306 508350
rect 417374 508294 417430 508350
rect 417498 508294 417554 508350
rect 417622 508294 417678 508350
rect 417250 508170 417306 508226
rect 417374 508170 417430 508226
rect 417498 508170 417554 508226
rect 417622 508170 417678 508226
rect 417250 508046 417306 508102
rect 417374 508046 417430 508102
rect 417498 508046 417554 508102
rect 417622 508046 417678 508102
rect 417250 507922 417306 507978
rect 417374 507922 417430 507978
rect 417498 507922 417554 507978
rect 417622 507922 417678 507978
rect 417250 490294 417306 490350
rect 417374 490294 417430 490350
rect 417498 490294 417554 490350
rect 417622 490294 417678 490350
rect 417250 490170 417306 490226
rect 417374 490170 417430 490226
rect 417498 490170 417554 490226
rect 417622 490170 417678 490226
rect 417250 490046 417306 490102
rect 417374 490046 417430 490102
rect 417498 490046 417554 490102
rect 417622 490046 417678 490102
rect 417250 489922 417306 489978
rect 417374 489922 417430 489978
rect 417498 489922 417554 489978
rect 417622 489922 417678 489978
rect 417250 472294 417306 472350
rect 417374 472294 417430 472350
rect 417498 472294 417554 472350
rect 417622 472294 417678 472350
rect 417250 472170 417306 472226
rect 417374 472170 417430 472226
rect 417498 472170 417554 472226
rect 417622 472170 417678 472226
rect 417250 472046 417306 472102
rect 417374 472046 417430 472102
rect 417498 472046 417554 472102
rect 417622 472046 417678 472102
rect 417250 471922 417306 471978
rect 417374 471922 417430 471978
rect 417498 471922 417554 471978
rect 417622 471922 417678 471978
rect 417250 454294 417306 454350
rect 417374 454294 417430 454350
rect 417498 454294 417554 454350
rect 417622 454294 417678 454350
rect 417250 454170 417306 454226
rect 417374 454170 417430 454226
rect 417498 454170 417554 454226
rect 417622 454170 417678 454226
rect 417250 454046 417306 454102
rect 417374 454046 417430 454102
rect 417498 454046 417554 454102
rect 417622 454046 417678 454102
rect 417250 453922 417306 453978
rect 417374 453922 417430 453978
rect 417498 453922 417554 453978
rect 417622 453922 417678 453978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 420970 514294 421026 514350
rect 421094 514294 421150 514350
rect 421218 514294 421274 514350
rect 421342 514294 421398 514350
rect 420970 514170 421026 514226
rect 421094 514170 421150 514226
rect 421218 514170 421274 514226
rect 421342 514170 421398 514226
rect 420970 514046 421026 514102
rect 421094 514046 421150 514102
rect 421218 514046 421274 514102
rect 421342 514046 421398 514102
rect 420970 513922 421026 513978
rect 421094 513922 421150 513978
rect 421218 513922 421274 513978
rect 421342 513922 421398 513978
rect 420970 496294 421026 496350
rect 421094 496294 421150 496350
rect 421218 496294 421274 496350
rect 421342 496294 421398 496350
rect 420970 496170 421026 496226
rect 421094 496170 421150 496226
rect 421218 496170 421274 496226
rect 421342 496170 421398 496226
rect 420970 496046 421026 496102
rect 421094 496046 421150 496102
rect 421218 496046 421274 496102
rect 421342 496046 421398 496102
rect 420970 495922 421026 495978
rect 421094 495922 421150 495978
rect 421218 495922 421274 495978
rect 421342 495922 421398 495978
rect 420970 478294 421026 478350
rect 421094 478294 421150 478350
rect 421218 478294 421274 478350
rect 421342 478294 421398 478350
rect 420970 478170 421026 478226
rect 421094 478170 421150 478226
rect 421218 478170 421274 478226
rect 421342 478170 421398 478226
rect 420970 478046 421026 478102
rect 421094 478046 421150 478102
rect 421218 478046 421274 478102
rect 421342 478046 421398 478102
rect 420970 477922 421026 477978
rect 421094 477922 421150 477978
rect 421218 477922 421274 477978
rect 421342 477922 421398 477978
rect 420970 460294 421026 460350
rect 421094 460294 421150 460350
rect 421218 460294 421274 460350
rect 421342 460294 421398 460350
rect 420970 460170 421026 460226
rect 421094 460170 421150 460226
rect 421218 460170 421274 460226
rect 421342 460170 421398 460226
rect 420970 460046 421026 460102
rect 421094 460046 421150 460102
rect 421218 460046 421274 460102
rect 421342 460046 421398 460102
rect 420970 459922 421026 459978
rect 421094 459922 421150 459978
rect 421218 459922 421274 459978
rect 421342 459922 421398 459978
rect 420970 442294 421026 442350
rect 421094 442294 421150 442350
rect 421218 442294 421274 442350
rect 421342 442294 421398 442350
rect 420970 442170 421026 442226
rect 421094 442170 421150 442226
rect 421218 442170 421274 442226
rect 421342 442170 421398 442226
rect 420970 442046 421026 442102
rect 421094 442046 421150 442102
rect 421218 442046 421274 442102
rect 421342 442046 421398 442102
rect 420970 441922 421026 441978
rect 421094 441922 421150 441978
rect 421218 441922 421274 441978
rect 421342 441922 421398 441978
rect 402970 424294 403026 424350
rect 403094 424294 403150 424350
rect 403218 424294 403274 424350
rect 403342 424294 403398 424350
rect 402970 424170 403026 424226
rect 403094 424170 403150 424226
rect 403218 424170 403274 424226
rect 403342 424170 403398 424226
rect 402970 424046 403026 424102
rect 403094 424046 403150 424102
rect 403218 424046 403274 424102
rect 403342 424046 403398 424102
rect 402970 423922 403026 423978
rect 403094 423922 403150 423978
rect 403218 423922 403274 423978
rect 403342 423922 403398 423978
rect 399250 418294 399306 418350
rect 399374 418294 399430 418350
rect 399498 418294 399554 418350
rect 399622 418294 399678 418350
rect 399250 418170 399306 418226
rect 399374 418170 399430 418226
rect 399498 418170 399554 418226
rect 399622 418170 399678 418226
rect 399250 418046 399306 418102
rect 399374 418046 399430 418102
rect 399498 418046 399554 418102
rect 399622 418046 399678 418102
rect 399250 417922 399306 417978
rect 399374 417922 399430 417978
rect 399498 417922 399554 417978
rect 399622 417922 399678 417978
rect 384970 406294 385026 406350
rect 385094 406294 385150 406350
rect 385218 406294 385274 406350
rect 385342 406294 385398 406350
rect 384970 406170 385026 406226
rect 385094 406170 385150 406226
rect 385218 406170 385274 406226
rect 385342 406170 385398 406226
rect 384970 406046 385026 406102
rect 385094 406046 385150 406102
rect 385218 406046 385274 406102
rect 385342 406046 385398 406102
rect 384970 405922 385026 405978
rect 385094 405922 385150 405978
rect 385218 405922 385274 405978
rect 385342 405922 385398 405978
rect 387078 406294 387134 406350
rect 387202 406294 387258 406350
rect 387078 406170 387134 406226
rect 387202 406170 387258 406226
rect 387078 406046 387134 406102
rect 387202 406046 387258 406102
rect 387078 405922 387134 405978
rect 387202 405922 387258 405978
rect 402438 418294 402494 418350
rect 402562 418294 402618 418350
rect 402438 418170 402494 418226
rect 402562 418170 402618 418226
rect 402438 418046 402494 418102
rect 402562 418046 402618 418102
rect 402438 417922 402494 417978
rect 402562 417922 402618 417978
rect 417798 424294 417854 424350
rect 417922 424294 417978 424350
rect 417798 424170 417854 424226
rect 417922 424170 417978 424226
rect 417798 424046 417854 424102
rect 417922 424046 417978 424102
rect 417798 423922 417854 423978
rect 417922 423922 417978 423978
rect 435250 597156 435306 597212
rect 435374 597156 435430 597212
rect 435498 597156 435554 597212
rect 435622 597156 435678 597212
rect 435250 597032 435306 597088
rect 435374 597032 435430 597088
rect 435498 597032 435554 597088
rect 435622 597032 435678 597088
rect 435250 596908 435306 596964
rect 435374 596908 435430 596964
rect 435498 596908 435554 596964
rect 435622 596908 435678 596964
rect 435250 596784 435306 596840
rect 435374 596784 435430 596840
rect 435498 596784 435554 596840
rect 435622 596784 435678 596840
rect 435250 580294 435306 580350
rect 435374 580294 435430 580350
rect 435498 580294 435554 580350
rect 435622 580294 435678 580350
rect 435250 580170 435306 580226
rect 435374 580170 435430 580226
rect 435498 580170 435554 580226
rect 435622 580170 435678 580226
rect 435250 580046 435306 580102
rect 435374 580046 435430 580102
rect 435498 580046 435554 580102
rect 435622 580046 435678 580102
rect 435250 579922 435306 579978
rect 435374 579922 435430 579978
rect 435498 579922 435554 579978
rect 435622 579922 435678 579978
rect 435250 562294 435306 562350
rect 435374 562294 435430 562350
rect 435498 562294 435554 562350
rect 435622 562294 435678 562350
rect 435250 562170 435306 562226
rect 435374 562170 435430 562226
rect 435498 562170 435554 562226
rect 435622 562170 435678 562226
rect 435250 562046 435306 562102
rect 435374 562046 435430 562102
rect 435498 562046 435554 562102
rect 435622 562046 435678 562102
rect 435250 561922 435306 561978
rect 435374 561922 435430 561978
rect 435498 561922 435554 561978
rect 435622 561922 435678 561978
rect 435250 544294 435306 544350
rect 435374 544294 435430 544350
rect 435498 544294 435554 544350
rect 435622 544294 435678 544350
rect 435250 544170 435306 544226
rect 435374 544170 435430 544226
rect 435498 544170 435554 544226
rect 435622 544170 435678 544226
rect 435250 544046 435306 544102
rect 435374 544046 435430 544102
rect 435498 544046 435554 544102
rect 435622 544046 435678 544102
rect 435250 543922 435306 543978
rect 435374 543922 435430 543978
rect 435498 543922 435554 543978
rect 435622 543922 435678 543978
rect 435250 526294 435306 526350
rect 435374 526294 435430 526350
rect 435498 526294 435554 526350
rect 435622 526294 435678 526350
rect 435250 526170 435306 526226
rect 435374 526170 435430 526226
rect 435498 526170 435554 526226
rect 435622 526170 435678 526226
rect 435250 526046 435306 526102
rect 435374 526046 435430 526102
rect 435498 526046 435554 526102
rect 435622 526046 435678 526102
rect 435250 525922 435306 525978
rect 435374 525922 435430 525978
rect 435498 525922 435554 525978
rect 435622 525922 435678 525978
rect 435250 508294 435306 508350
rect 435374 508294 435430 508350
rect 435498 508294 435554 508350
rect 435622 508294 435678 508350
rect 435250 508170 435306 508226
rect 435374 508170 435430 508226
rect 435498 508170 435554 508226
rect 435622 508170 435678 508226
rect 435250 508046 435306 508102
rect 435374 508046 435430 508102
rect 435498 508046 435554 508102
rect 435622 508046 435678 508102
rect 435250 507922 435306 507978
rect 435374 507922 435430 507978
rect 435498 507922 435554 507978
rect 435622 507922 435678 507978
rect 435250 490294 435306 490350
rect 435374 490294 435430 490350
rect 435498 490294 435554 490350
rect 435622 490294 435678 490350
rect 435250 490170 435306 490226
rect 435374 490170 435430 490226
rect 435498 490170 435554 490226
rect 435622 490170 435678 490226
rect 435250 490046 435306 490102
rect 435374 490046 435430 490102
rect 435498 490046 435554 490102
rect 435622 490046 435678 490102
rect 435250 489922 435306 489978
rect 435374 489922 435430 489978
rect 435498 489922 435554 489978
rect 435622 489922 435678 489978
rect 435250 472294 435306 472350
rect 435374 472294 435430 472350
rect 435498 472294 435554 472350
rect 435622 472294 435678 472350
rect 435250 472170 435306 472226
rect 435374 472170 435430 472226
rect 435498 472170 435554 472226
rect 435622 472170 435678 472226
rect 435250 472046 435306 472102
rect 435374 472046 435430 472102
rect 435498 472046 435554 472102
rect 435622 472046 435678 472102
rect 435250 471922 435306 471978
rect 435374 471922 435430 471978
rect 435498 471922 435554 471978
rect 435622 471922 435678 471978
rect 435250 454294 435306 454350
rect 435374 454294 435430 454350
rect 435498 454294 435554 454350
rect 435622 454294 435678 454350
rect 435250 454170 435306 454226
rect 435374 454170 435430 454226
rect 435498 454170 435554 454226
rect 435622 454170 435678 454226
rect 435250 454046 435306 454102
rect 435374 454046 435430 454102
rect 435498 454046 435554 454102
rect 435622 454046 435678 454102
rect 435250 453922 435306 453978
rect 435374 453922 435430 453978
rect 435498 453922 435554 453978
rect 435622 453922 435678 453978
rect 433158 436261 433214 436317
rect 433282 436261 433338 436317
rect 433158 436137 433214 436193
rect 433282 436137 433338 436193
rect 433158 436013 433214 436069
rect 433282 436013 433338 436069
rect 433158 435889 433214 435945
rect 433282 435889 433338 435945
rect 435250 436294 435306 436350
rect 435374 436294 435430 436350
rect 435498 436294 435554 436350
rect 435622 436294 435678 436350
rect 435250 436170 435306 436226
rect 435374 436170 435430 436226
rect 435498 436170 435554 436226
rect 435622 436170 435678 436226
rect 435250 436046 435306 436102
rect 435374 436046 435430 436102
rect 435498 436046 435554 436102
rect 435622 436046 435678 436102
rect 435250 435922 435306 435978
rect 435374 435922 435430 435978
rect 435498 435922 435554 435978
rect 435622 435922 435678 435978
rect 420970 424294 421026 424350
rect 421094 424294 421150 424350
rect 421218 424294 421274 424350
rect 421342 424294 421398 424350
rect 420970 424170 421026 424226
rect 421094 424170 421150 424226
rect 421218 424170 421274 424226
rect 421342 424170 421398 424226
rect 420970 424046 421026 424102
rect 421094 424046 421150 424102
rect 421218 424046 421274 424102
rect 421342 424046 421398 424102
rect 420970 423922 421026 423978
rect 421094 423922 421150 423978
rect 421218 423922 421274 423978
rect 421342 423922 421398 423978
rect 402970 406294 403026 406350
rect 403094 406294 403150 406350
rect 403218 406294 403274 406350
rect 403342 406294 403398 406350
rect 402970 406170 403026 406226
rect 403094 406170 403150 406226
rect 403218 406170 403274 406226
rect 403342 406170 403398 406226
rect 402970 406046 403026 406102
rect 403094 406046 403150 406102
rect 403218 406046 403274 406102
rect 403342 406046 403398 406102
rect 402970 405922 403026 405978
rect 403094 405922 403150 405978
rect 403218 405922 403274 405978
rect 403342 405922 403398 405978
rect 399250 400294 399306 400350
rect 399374 400294 399430 400350
rect 399498 400294 399554 400350
rect 399622 400294 399678 400350
rect 399250 400170 399306 400226
rect 399374 400170 399430 400226
rect 399498 400170 399554 400226
rect 399622 400170 399678 400226
rect 399250 400046 399306 400102
rect 399374 400046 399430 400102
rect 399498 400046 399554 400102
rect 399622 400046 399678 400102
rect 399250 399922 399306 399978
rect 399374 399922 399430 399978
rect 399498 399922 399554 399978
rect 399622 399922 399678 399978
rect 384970 388294 385026 388350
rect 385094 388294 385150 388350
rect 385218 388294 385274 388350
rect 385342 388294 385398 388350
rect 384970 388170 385026 388226
rect 385094 388170 385150 388226
rect 385218 388170 385274 388226
rect 385342 388170 385398 388226
rect 384970 388046 385026 388102
rect 385094 388046 385150 388102
rect 385218 388046 385274 388102
rect 385342 388046 385398 388102
rect 384970 387922 385026 387978
rect 385094 387922 385150 387978
rect 385218 387922 385274 387978
rect 385342 387922 385398 387978
rect 387078 388294 387134 388350
rect 387202 388294 387258 388350
rect 387078 388170 387134 388226
rect 387202 388170 387258 388226
rect 387078 388046 387134 388102
rect 387202 388046 387258 388102
rect 387078 387922 387134 387978
rect 387202 387922 387258 387978
rect 402438 400294 402494 400350
rect 402562 400294 402618 400350
rect 402438 400170 402494 400226
rect 402562 400170 402618 400226
rect 402438 400046 402494 400102
rect 402562 400046 402618 400102
rect 402438 399922 402494 399978
rect 402562 399922 402618 399978
rect 417798 406294 417854 406350
rect 417922 406294 417978 406350
rect 417798 406170 417854 406226
rect 417922 406170 417978 406226
rect 417798 406046 417854 406102
rect 417922 406046 417978 406102
rect 417798 405922 417854 405978
rect 417922 405922 417978 405978
rect 433158 418294 433214 418350
rect 433282 418294 433338 418350
rect 433158 418170 433214 418226
rect 433282 418170 433338 418226
rect 433158 418046 433214 418102
rect 433282 418046 433338 418102
rect 433158 417922 433214 417978
rect 433282 417922 433338 417978
rect 435250 418294 435306 418350
rect 435374 418294 435430 418350
rect 435498 418294 435554 418350
rect 435622 418294 435678 418350
rect 435250 418170 435306 418226
rect 435374 418170 435430 418226
rect 435498 418170 435554 418226
rect 435622 418170 435678 418226
rect 435250 418046 435306 418102
rect 435374 418046 435430 418102
rect 435498 418046 435554 418102
rect 435622 418046 435678 418102
rect 435250 417922 435306 417978
rect 435374 417922 435430 417978
rect 435498 417922 435554 417978
rect 435622 417922 435678 417978
rect 420970 406294 421026 406350
rect 421094 406294 421150 406350
rect 421218 406294 421274 406350
rect 421342 406294 421398 406350
rect 420970 406170 421026 406226
rect 421094 406170 421150 406226
rect 421218 406170 421274 406226
rect 421342 406170 421398 406226
rect 420970 406046 421026 406102
rect 421094 406046 421150 406102
rect 421218 406046 421274 406102
rect 421342 406046 421398 406102
rect 420970 405922 421026 405978
rect 421094 405922 421150 405978
rect 421218 405922 421274 405978
rect 421342 405922 421398 405978
rect 402970 388294 403026 388350
rect 403094 388294 403150 388350
rect 403218 388294 403274 388350
rect 403342 388294 403398 388350
rect 402970 388170 403026 388226
rect 403094 388170 403150 388226
rect 403218 388170 403274 388226
rect 403342 388170 403398 388226
rect 402970 388046 403026 388102
rect 403094 388046 403150 388102
rect 403218 388046 403274 388102
rect 403342 388046 403398 388102
rect 402970 387922 403026 387978
rect 403094 387922 403150 387978
rect 403218 387922 403274 387978
rect 403342 387922 403398 387978
rect 399250 382294 399306 382350
rect 399374 382294 399430 382350
rect 399498 382294 399554 382350
rect 399622 382294 399678 382350
rect 399250 382170 399306 382226
rect 399374 382170 399430 382226
rect 399498 382170 399554 382226
rect 399622 382170 399678 382226
rect 399250 382046 399306 382102
rect 399374 382046 399430 382102
rect 399498 382046 399554 382102
rect 399622 382046 399678 382102
rect 399250 381922 399306 381978
rect 399374 381922 399430 381978
rect 399498 381922 399554 381978
rect 399622 381922 399678 381978
rect 384970 370294 385026 370350
rect 385094 370294 385150 370350
rect 385218 370294 385274 370350
rect 385342 370294 385398 370350
rect 384970 370170 385026 370226
rect 385094 370170 385150 370226
rect 385218 370170 385274 370226
rect 385342 370170 385398 370226
rect 384970 370046 385026 370102
rect 385094 370046 385150 370102
rect 385218 370046 385274 370102
rect 385342 370046 385398 370102
rect 384970 369922 385026 369978
rect 385094 369922 385150 369978
rect 385218 369922 385274 369978
rect 385342 369922 385398 369978
rect 387078 370294 387134 370350
rect 387202 370294 387258 370350
rect 387078 370170 387134 370226
rect 387202 370170 387258 370226
rect 387078 370046 387134 370102
rect 387202 370046 387258 370102
rect 387078 369922 387134 369978
rect 387202 369922 387258 369978
rect 402438 382294 402494 382350
rect 402562 382294 402618 382350
rect 402438 382170 402494 382226
rect 402562 382170 402618 382226
rect 402438 382046 402494 382102
rect 402562 382046 402618 382102
rect 402438 381922 402494 381978
rect 402562 381922 402618 381978
rect 417798 388294 417854 388350
rect 417922 388294 417978 388350
rect 417798 388170 417854 388226
rect 417922 388170 417978 388226
rect 417798 388046 417854 388102
rect 417922 388046 417978 388102
rect 417798 387922 417854 387978
rect 417922 387922 417978 387978
rect 433158 400294 433214 400350
rect 433282 400294 433338 400350
rect 433158 400170 433214 400226
rect 433282 400170 433338 400226
rect 433158 400046 433214 400102
rect 433282 400046 433338 400102
rect 433158 399922 433214 399978
rect 433282 399922 433338 399978
rect 435250 400294 435306 400350
rect 435374 400294 435430 400350
rect 435498 400294 435554 400350
rect 435622 400294 435678 400350
rect 435250 400170 435306 400226
rect 435374 400170 435430 400226
rect 435498 400170 435554 400226
rect 435622 400170 435678 400226
rect 435250 400046 435306 400102
rect 435374 400046 435430 400102
rect 435498 400046 435554 400102
rect 435622 400046 435678 400102
rect 435250 399922 435306 399978
rect 435374 399922 435430 399978
rect 435498 399922 435554 399978
rect 435622 399922 435678 399978
rect 420970 388294 421026 388350
rect 421094 388294 421150 388350
rect 421218 388294 421274 388350
rect 421342 388294 421398 388350
rect 420970 388170 421026 388226
rect 421094 388170 421150 388226
rect 421218 388170 421274 388226
rect 421342 388170 421398 388226
rect 420970 388046 421026 388102
rect 421094 388046 421150 388102
rect 421218 388046 421274 388102
rect 421342 388046 421398 388102
rect 420970 387922 421026 387978
rect 421094 387922 421150 387978
rect 421218 387922 421274 387978
rect 421342 387922 421398 387978
rect 402970 370294 403026 370350
rect 403094 370294 403150 370350
rect 403218 370294 403274 370350
rect 403342 370294 403398 370350
rect 402970 370170 403026 370226
rect 403094 370170 403150 370226
rect 403218 370170 403274 370226
rect 403342 370170 403398 370226
rect 402970 370046 403026 370102
rect 403094 370046 403150 370102
rect 403218 370046 403274 370102
rect 403342 370046 403398 370102
rect 402970 369922 403026 369978
rect 403094 369922 403150 369978
rect 403218 369922 403274 369978
rect 403342 369922 403398 369978
rect 399250 364294 399306 364350
rect 399374 364294 399430 364350
rect 399498 364294 399554 364350
rect 399622 364294 399678 364350
rect 399250 364170 399306 364226
rect 399374 364170 399430 364226
rect 399498 364170 399554 364226
rect 399622 364170 399678 364226
rect 399250 364046 399306 364102
rect 399374 364046 399430 364102
rect 399498 364046 399554 364102
rect 399622 364046 399678 364102
rect 399250 363922 399306 363978
rect 399374 363922 399430 363978
rect 399498 363922 399554 363978
rect 399622 363922 399678 363978
rect 384970 352294 385026 352350
rect 385094 352294 385150 352350
rect 385218 352294 385274 352350
rect 385342 352294 385398 352350
rect 384970 352170 385026 352226
rect 385094 352170 385150 352226
rect 385218 352170 385274 352226
rect 385342 352170 385398 352226
rect 384970 352046 385026 352102
rect 385094 352046 385150 352102
rect 385218 352046 385274 352102
rect 385342 352046 385398 352102
rect 384970 351922 385026 351978
rect 385094 351922 385150 351978
rect 385218 351922 385274 351978
rect 385342 351922 385398 351978
rect 387078 352294 387134 352350
rect 387202 352294 387258 352350
rect 387078 352170 387134 352226
rect 387202 352170 387258 352226
rect 387078 352046 387134 352102
rect 387202 352046 387258 352102
rect 387078 351922 387134 351978
rect 387202 351922 387258 351978
rect 402438 364294 402494 364350
rect 402562 364294 402618 364350
rect 402438 364170 402494 364226
rect 402562 364170 402618 364226
rect 402438 364046 402494 364102
rect 402562 364046 402618 364102
rect 402438 363922 402494 363978
rect 402562 363922 402618 363978
rect 417798 370294 417854 370350
rect 417922 370294 417978 370350
rect 417798 370170 417854 370226
rect 417922 370170 417978 370226
rect 417798 370046 417854 370102
rect 417922 370046 417978 370102
rect 417798 369922 417854 369978
rect 417922 369922 417978 369978
rect 433158 382294 433214 382350
rect 433282 382294 433338 382350
rect 433158 382170 433214 382226
rect 433282 382170 433338 382226
rect 433158 382046 433214 382102
rect 433282 382046 433338 382102
rect 433158 381922 433214 381978
rect 433282 381922 433338 381978
rect 435250 382294 435306 382350
rect 435374 382294 435430 382350
rect 435498 382294 435554 382350
rect 435622 382294 435678 382350
rect 435250 382170 435306 382226
rect 435374 382170 435430 382226
rect 435498 382170 435554 382226
rect 435622 382170 435678 382226
rect 435250 382046 435306 382102
rect 435374 382046 435430 382102
rect 435498 382046 435554 382102
rect 435622 382046 435678 382102
rect 435250 381922 435306 381978
rect 435374 381922 435430 381978
rect 435498 381922 435554 381978
rect 435622 381922 435678 381978
rect 420970 370294 421026 370350
rect 421094 370294 421150 370350
rect 421218 370294 421274 370350
rect 421342 370294 421398 370350
rect 420970 370170 421026 370226
rect 421094 370170 421150 370226
rect 421218 370170 421274 370226
rect 421342 370170 421398 370226
rect 420970 370046 421026 370102
rect 421094 370046 421150 370102
rect 421218 370046 421274 370102
rect 421342 370046 421398 370102
rect 420970 369922 421026 369978
rect 421094 369922 421150 369978
rect 421218 369922 421274 369978
rect 421342 369922 421398 369978
rect 402970 352294 403026 352350
rect 403094 352294 403150 352350
rect 403218 352294 403274 352350
rect 403342 352294 403398 352350
rect 402970 352170 403026 352226
rect 403094 352170 403150 352226
rect 403218 352170 403274 352226
rect 403342 352170 403398 352226
rect 402970 352046 403026 352102
rect 403094 352046 403150 352102
rect 403218 352046 403274 352102
rect 403342 352046 403398 352102
rect 402970 351922 403026 351978
rect 403094 351922 403150 351978
rect 403218 351922 403274 351978
rect 403342 351922 403398 351978
rect 399250 346294 399306 346350
rect 399374 346294 399430 346350
rect 399498 346294 399554 346350
rect 399622 346294 399678 346350
rect 399250 346170 399306 346226
rect 399374 346170 399430 346226
rect 399498 346170 399554 346226
rect 399622 346170 399678 346226
rect 399250 346046 399306 346102
rect 399374 346046 399430 346102
rect 399498 346046 399554 346102
rect 399622 346046 399678 346102
rect 399250 345922 399306 345978
rect 399374 345922 399430 345978
rect 399498 345922 399554 345978
rect 399622 345922 399678 345978
rect 384970 334294 385026 334350
rect 385094 334294 385150 334350
rect 385218 334294 385274 334350
rect 385342 334294 385398 334350
rect 384970 334170 385026 334226
rect 385094 334170 385150 334226
rect 385218 334170 385274 334226
rect 385342 334170 385398 334226
rect 384970 334046 385026 334102
rect 385094 334046 385150 334102
rect 385218 334046 385274 334102
rect 385342 334046 385398 334102
rect 384970 333922 385026 333978
rect 385094 333922 385150 333978
rect 385218 333922 385274 333978
rect 385342 333922 385398 333978
rect 387078 334294 387134 334350
rect 387202 334294 387258 334350
rect 387078 334170 387134 334226
rect 387202 334170 387258 334226
rect 387078 334046 387134 334102
rect 387202 334046 387258 334102
rect 387078 333922 387134 333978
rect 387202 333922 387258 333978
rect 402438 346294 402494 346350
rect 402562 346294 402618 346350
rect 402438 346170 402494 346226
rect 402562 346170 402618 346226
rect 402438 346046 402494 346102
rect 402562 346046 402618 346102
rect 402438 345922 402494 345978
rect 402562 345922 402618 345978
rect 417798 352294 417854 352350
rect 417922 352294 417978 352350
rect 417798 352170 417854 352226
rect 417922 352170 417978 352226
rect 417798 352046 417854 352102
rect 417922 352046 417978 352102
rect 417798 351922 417854 351978
rect 417922 351922 417978 351978
rect 433158 364294 433214 364350
rect 433282 364294 433338 364350
rect 433158 364170 433214 364226
rect 433282 364170 433338 364226
rect 433158 364046 433214 364102
rect 433282 364046 433338 364102
rect 433158 363922 433214 363978
rect 433282 363922 433338 363978
rect 435250 364294 435306 364350
rect 435374 364294 435430 364350
rect 435498 364294 435554 364350
rect 435622 364294 435678 364350
rect 435250 364170 435306 364226
rect 435374 364170 435430 364226
rect 435498 364170 435554 364226
rect 435622 364170 435678 364226
rect 435250 364046 435306 364102
rect 435374 364046 435430 364102
rect 435498 364046 435554 364102
rect 435622 364046 435678 364102
rect 435250 363922 435306 363978
rect 435374 363922 435430 363978
rect 435498 363922 435554 363978
rect 435622 363922 435678 363978
rect 420970 352294 421026 352350
rect 421094 352294 421150 352350
rect 421218 352294 421274 352350
rect 421342 352294 421398 352350
rect 420970 352170 421026 352226
rect 421094 352170 421150 352226
rect 421218 352170 421274 352226
rect 421342 352170 421398 352226
rect 420970 352046 421026 352102
rect 421094 352046 421150 352102
rect 421218 352046 421274 352102
rect 421342 352046 421398 352102
rect 420970 351922 421026 351978
rect 421094 351922 421150 351978
rect 421218 351922 421274 351978
rect 421342 351922 421398 351978
rect 402970 334294 403026 334350
rect 403094 334294 403150 334350
rect 403218 334294 403274 334350
rect 403342 334294 403398 334350
rect 402970 334170 403026 334226
rect 403094 334170 403150 334226
rect 403218 334170 403274 334226
rect 403342 334170 403398 334226
rect 402970 334046 403026 334102
rect 403094 334046 403150 334102
rect 403218 334046 403274 334102
rect 403342 334046 403398 334102
rect 402970 333922 403026 333978
rect 403094 333922 403150 333978
rect 403218 333922 403274 333978
rect 403342 333922 403398 333978
rect 399250 328294 399306 328350
rect 399374 328294 399430 328350
rect 399498 328294 399554 328350
rect 399622 328294 399678 328350
rect 399250 328170 399306 328226
rect 399374 328170 399430 328226
rect 399498 328170 399554 328226
rect 399622 328170 399678 328226
rect 399250 328046 399306 328102
rect 399374 328046 399430 328102
rect 399498 328046 399554 328102
rect 399622 328046 399678 328102
rect 399250 327922 399306 327978
rect 399374 327922 399430 327978
rect 399498 327922 399554 327978
rect 399622 327922 399678 327978
rect 384970 316294 385026 316350
rect 385094 316294 385150 316350
rect 385218 316294 385274 316350
rect 385342 316294 385398 316350
rect 384970 316170 385026 316226
rect 385094 316170 385150 316226
rect 385218 316170 385274 316226
rect 385342 316170 385398 316226
rect 384970 316046 385026 316102
rect 385094 316046 385150 316102
rect 385218 316046 385274 316102
rect 385342 316046 385398 316102
rect 384970 315922 385026 315978
rect 385094 315922 385150 315978
rect 385218 315922 385274 315978
rect 385342 315922 385398 315978
rect 387078 316294 387134 316350
rect 387202 316294 387258 316350
rect 387078 316170 387134 316226
rect 387202 316170 387258 316226
rect 387078 316046 387134 316102
rect 387202 316046 387258 316102
rect 387078 315922 387134 315978
rect 387202 315922 387258 315978
rect 402438 328294 402494 328350
rect 402562 328294 402618 328350
rect 402438 328170 402494 328226
rect 402562 328170 402618 328226
rect 402438 328046 402494 328102
rect 402562 328046 402618 328102
rect 402438 327922 402494 327978
rect 402562 327922 402618 327978
rect 417798 334294 417854 334350
rect 417922 334294 417978 334350
rect 417798 334170 417854 334226
rect 417922 334170 417978 334226
rect 417798 334046 417854 334102
rect 417922 334046 417978 334102
rect 417798 333922 417854 333978
rect 417922 333922 417978 333978
rect 433158 346294 433214 346350
rect 433282 346294 433338 346350
rect 433158 346170 433214 346226
rect 433282 346170 433338 346226
rect 433158 346046 433214 346102
rect 433282 346046 433338 346102
rect 433158 345922 433214 345978
rect 433282 345922 433338 345978
rect 435250 346294 435306 346350
rect 435374 346294 435430 346350
rect 435498 346294 435554 346350
rect 435622 346294 435678 346350
rect 435250 346170 435306 346226
rect 435374 346170 435430 346226
rect 435498 346170 435554 346226
rect 435622 346170 435678 346226
rect 435250 346046 435306 346102
rect 435374 346046 435430 346102
rect 435498 346046 435554 346102
rect 435622 346046 435678 346102
rect 435250 345922 435306 345978
rect 435374 345922 435430 345978
rect 435498 345922 435554 345978
rect 435622 345922 435678 345978
rect 420970 334294 421026 334350
rect 421094 334294 421150 334350
rect 421218 334294 421274 334350
rect 421342 334294 421398 334350
rect 420970 334170 421026 334226
rect 421094 334170 421150 334226
rect 421218 334170 421274 334226
rect 421342 334170 421398 334226
rect 420970 334046 421026 334102
rect 421094 334046 421150 334102
rect 421218 334046 421274 334102
rect 421342 334046 421398 334102
rect 420970 333922 421026 333978
rect 421094 333922 421150 333978
rect 421218 333922 421274 333978
rect 421342 333922 421398 333978
rect 402970 316294 403026 316350
rect 403094 316294 403150 316350
rect 403218 316294 403274 316350
rect 403342 316294 403398 316350
rect 402970 316170 403026 316226
rect 403094 316170 403150 316226
rect 403218 316170 403274 316226
rect 403342 316170 403398 316226
rect 402970 316046 403026 316102
rect 403094 316046 403150 316102
rect 403218 316046 403274 316102
rect 403342 316046 403398 316102
rect 402970 315922 403026 315978
rect 403094 315922 403150 315978
rect 403218 315922 403274 315978
rect 403342 315922 403398 315978
rect 399250 310294 399306 310350
rect 399374 310294 399430 310350
rect 399498 310294 399554 310350
rect 399622 310294 399678 310350
rect 399250 310170 399306 310226
rect 399374 310170 399430 310226
rect 399498 310170 399554 310226
rect 399622 310170 399678 310226
rect 399250 310046 399306 310102
rect 399374 310046 399430 310102
rect 399498 310046 399554 310102
rect 399622 310046 399678 310102
rect 399250 309922 399306 309978
rect 399374 309922 399430 309978
rect 399498 309922 399554 309978
rect 399622 309922 399678 309978
rect 384970 298294 385026 298350
rect 385094 298294 385150 298350
rect 385218 298294 385274 298350
rect 385342 298294 385398 298350
rect 384970 298170 385026 298226
rect 385094 298170 385150 298226
rect 385218 298170 385274 298226
rect 385342 298170 385398 298226
rect 384970 298046 385026 298102
rect 385094 298046 385150 298102
rect 385218 298046 385274 298102
rect 385342 298046 385398 298102
rect 384970 297922 385026 297978
rect 385094 297922 385150 297978
rect 385218 297922 385274 297978
rect 385342 297922 385398 297978
rect 387078 298294 387134 298350
rect 387202 298294 387258 298350
rect 387078 298170 387134 298226
rect 387202 298170 387258 298226
rect 387078 298046 387134 298102
rect 387202 298046 387258 298102
rect 387078 297922 387134 297978
rect 387202 297922 387258 297978
rect 402438 310294 402494 310350
rect 402562 310294 402618 310350
rect 402438 310170 402494 310226
rect 402562 310170 402618 310226
rect 402438 310046 402494 310102
rect 402562 310046 402618 310102
rect 402438 309922 402494 309978
rect 402562 309922 402618 309978
rect 417798 316294 417854 316350
rect 417922 316294 417978 316350
rect 417798 316170 417854 316226
rect 417922 316170 417978 316226
rect 417798 316046 417854 316102
rect 417922 316046 417978 316102
rect 417798 315922 417854 315978
rect 417922 315922 417978 315978
rect 433158 328294 433214 328350
rect 433282 328294 433338 328350
rect 433158 328170 433214 328226
rect 433282 328170 433338 328226
rect 433158 328046 433214 328102
rect 433282 328046 433338 328102
rect 433158 327922 433214 327978
rect 433282 327922 433338 327978
rect 435250 328294 435306 328350
rect 435374 328294 435430 328350
rect 435498 328294 435554 328350
rect 435622 328294 435678 328350
rect 435250 328170 435306 328226
rect 435374 328170 435430 328226
rect 435498 328170 435554 328226
rect 435622 328170 435678 328226
rect 435250 328046 435306 328102
rect 435374 328046 435430 328102
rect 435498 328046 435554 328102
rect 435622 328046 435678 328102
rect 435250 327922 435306 327978
rect 435374 327922 435430 327978
rect 435498 327922 435554 327978
rect 435622 327922 435678 327978
rect 420970 316294 421026 316350
rect 421094 316294 421150 316350
rect 421218 316294 421274 316350
rect 421342 316294 421398 316350
rect 420970 316170 421026 316226
rect 421094 316170 421150 316226
rect 421218 316170 421274 316226
rect 421342 316170 421398 316226
rect 420970 316046 421026 316102
rect 421094 316046 421150 316102
rect 421218 316046 421274 316102
rect 421342 316046 421398 316102
rect 420970 315922 421026 315978
rect 421094 315922 421150 315978
rect 421218 315922 421274 315978
rect 421342 315922 421398 315978
rect 402970 298294 403026 298350
rect 403094 298294 403150 298350
rect 403218 298294 403274 298350
rect 403342 298294 403398 298350
rect 402970 298170 403026 298226
rect 403094 298170 403150 298226
rect 403218 298170 403274 298226
rect 403342 298170 403398 298226
rect 402970 298046 403026 298102
rect 403094 298046 403150 298102
rect 403218 298046 403274 298102
rect 403342 298046 403398 298102
rect 402970 297922 403026 297978
rect 403094 297922 403150 297978
rect 403218 297922 403274 297978
rect 403342 297922 403398 297978
rect 399250 292294 399306 292350
rect 399374 292294 399430 292350
rect 399498 292294 399554 292350
rect 399622 292294 399678 292350
rect 399250 292170 399306 292226
rect 399374 292170 399430 292226
rect 399498 292170 399554 292226
rect 399622 292170 399678 292226
rect 399250 292046 399306 292102
rect 399374 292046 399430 292102
rect 399498 292046 399554 292102
rect 399622 292046 399678 292102
rect 399250 291922 399306 291978
rect 399374 291922 399430 291978
rect 399498 291922 399554 291978
rect 399622 291922 399678 291978
rect 384970 280294 385026 280350
rect 385094 280294 385150 280350
rect 385218 280294 385274 280350
rect 385342 280294 385398 280350
rect 384970 280170 385026 280226
rect 385094 280170 385150 280226
rect 385218 280170 385274 280226
rect 385342 280170 385398 280226
rect 384970 280046 385026 280102
rect 385094 280046 385150 280102
rect 385218 280046 385274 280102
rect 385342 280046 385398 280102
rect 384970 279922 385026 279978
rect 385094 279922 385150 279978
rect 385218 279922 385274 279978
rect 385342 279922 385398 279978
rect 387078 280294 387134 280350
rect 387202 280294 387258 280350
rect 387078 280170 387134 280226
rect 387202 280170 387258 280226
rect 387078 280046 387134 280102
rect 387202 280046 387258 280102
rect 387078 279922 387134 279978
rect 387202 279922 387258 279978
rect 402438 292294 402494 292350
rect 402562 292294 402618 292350
rect 402438 292170 402494 292226
rect 402562 292170 402618 292226
rect 402438 292046 402494 292102
rect 402562 292046 402618 292102
rect 402438 291922 402494 291978
rect 402562 291922 402618 291978
rect 417798 298294 417854 298350
rect 417922 298294 417978 298350
rect 417798 298170 417854 298226
rect 417922 298170 417978 298226
rect 417798 298046 417854 298102
rect 417922 298046 417978 298102
rect 417798 297922 417854 297978
rect 417922 297922 417978 297978
rect 433158 310294 433214 310350
rect 433282 310294 433338 310350
rect 433158 310170 433214 310226
rect 433282 310170 433338 310226
rect 433158 310046 433214 310102
rect 433282 310046 433338 310102
rect 433158 309922 433214 309978
rect 433282 309922 433338 309978
rect 435250 310294 435306 310350
rect 435374 310294 435430 310350
rect 435498 310294 435554 310350
rect 435622 310294 435678 310350
rect 435250 310170 435306 310226
rect 435374 310170 435430 310226
rect 435498 310170 435554 310226
rect 435622 310170 435678 310226
rect 435250 310046 435306 310102
rect 435374 310046 435430 310102
rect 435498 310046 435554 310102
rect 435622 310046 435678 310102
rect 435250 309922 435306 309978
rect 435374 309922 435430 309978
rect 435498 309922 435554 309978
rect 435622 309922 435678 309978
rect 420970 298294 421026 298350
rect 421094 298294 421150 298350
rect 421218 298294 421274 298350
rect 421342 298294 421398 298350
rect 420970 298170 421026 298226
rect 421094 298170 421150 298226
rect 421218 298170 421274 298226
rect 421342 298170 421398 298226
rect 420970 298046 421026 298102
rect 421094 298046 421150 298102
rect 421218 298046 421274 298102
rect 421342 298046 421398 298102
rect 420970 297922 421026 297978
rect 421094 297922 421150 297978
rect 421218 297922 421274 297978
rect 421342 297922 421398 297978
rect 402970 280294 403026 280350
rect 403094 280294 403150 280350
rect 403218 280294 403274 280350
rect 403342 280294 403398 280350
rect 402970 280170 403026 280226
rect 403094 280170 403150 280226
rect 403218 280170 403274 280226
rect 403342 280170 403398 280226
rect 402970 280046 403026 280102
rect 403094 280046 403150 280102
rect 403218 280046 403274 280102
rect 403342 280046 403398 280102
rect 402970 279922 403026 279978
rect 403094 279922 403150 279978
rect 403218 279922 403274 279978
rect 403342 279922 403398 279978
rect 399250 274294 399306 274350
rect 399374 274294 399430 274350
rect 399498 274294 399554 274350
rect 399622 274294 399678 274350
rect 399250 274170 399306 274226
rect 399374 274170 399430 274226
rect 399498 274170 399554 274226
rect 399622 274170 399678 274226
rect 399250 274046 399306 274102
rect 399374 274046 399430 274102
rect 399498 274046 399554 274102
rect 399622 274046 399678 274102
rect 399250 273922 399306 273978
rect 399374 273922 399430 273978
rect 399498 273922 399554 273978
rect 399622 273922 399678 273978
rect 384970 262294 385026 262350
rect 385094 262294 385150 262350
rect 385218 262294 385274 262350
rect 385342 262294 385398 262350
rect 384970 262170 385026 262226
rect 385094 262170 385150 262226
rect 385218 262170 385274 262226
rect 385342 262170 385398 262226
rect 384970 262046 385026 262102
rect 385094 262046 385150 262102
rect 385218 262046 385274 262102
rect 385342 262046 385398 262102
rect 384970 261922 385026 261978
rect 385094 261922 385150 261978
rect 385218 261922 385274 261978
rect 385342 261922 385398 261978
rect 387078 262294 387134 262350
rect 387202 262294 387258 262350
rect 387078 262170 387134 262226
rect 387202 262170 387258 262226
rect 387078 262046 387134 262102
rect 387202 262046 387258 262102
rect 387078 261922 387134 261978
rect 387202 261922 387258 261978
rect 402438 274294 402494 274350
rect 402562 274294 402618 274350
rect 402438 274170 402494 274226
rect 402562 274170 402618 274226
rect 402438 274046 402494 274102
rect 402562 274046 402618 274102
rect 402438 273922 402494 273978
rect 402562 273922 402618 273978
rect 417798 280294 417854 280350
rect 417922 280294 417978 280350
rect 417798 280170 417854 280226
rect 417922 280170 417978 280226
rect 417798 280046 417854 280102
rect 417922 280046 417978 280102
rect 417798 279922 417854 279978
rect 417922 279922 417978 279978
rect 433158 292294 433214 292350
rect 433282 292294 433338 292350
rect 433158 292170 433214 292226
rect 433282 292170 433338 292226
rect 433158 292046 433214 292102
rect 433282 292046 433338 292102
rect 433158 291922 433214 291978
rect 433282 291922 433338 291978
rect 435250 292294 435306 292350
rect 435374 292294 435430 292350
rect 435498 292294 435554 292350
rect 435622 292294 435678 292350
rect 435250 292170 435306 292226
rect 435374 292170 435430 292226
rect 435498 292170 435554 292226
rect 435622 292170 435678 292226
rect 435250 292046 435306 292102
rect 435374 292046 435430 292102
rect 435498 292046 435554 292102
rect 435622 292046 435678 292102
rect 435250 291922 435306 291978
rect 435374 291922 435430 291978
rect 435498 291922 435554 291978
rect 435622 291922 435678 291978
rect 420970 280294 421026 280350
rect 421094 280294 421150 280350
rect 421218 280294 421274 280350
rect 421342 280294 421398 280350
rect 420970 280170 421026 280226
rect 421094 280170 421150 280226
rect 421218 280170 421274 280226
rect 421342 280170 421398 280226
rect 420970 280046 421026 280102
rect 421094 280046 421150 280102
rect 421218 280046 421274 280102
rect 421342 280046 421398 280102
rect 420970 279922 421026 279978
rect 421094 279922 421150 279978
rect 421218 279922 421274 279978
rect 421342 279922 421398 279978
rect 402970 262294 403026 262350
rect 403094 262294 403150 262350
rect 403218 262294 403274 262350
rect 403342 262294 403398 262350
rect 402970 262170 403026 262226
rect 403094 262170 403150 262226
rect 403218 262170 403274 262226
rect 403342 262170 403398 262226
rect 402970 262046 403026 262102
rect 403094 262046 403150 262102
rect 403218 262046 403274 262102
rect 403342 262046 403398 262102
rect 402970 261922 403026 261978
rect 403094 261922 403150 261978
rect 403218 261922 403274 261978
rect 403342 261922 403398 261978
rect 399250 256294 399306 256350
rect 399374 256294 399430 256350
rect 399498 256294 399554 256350
rect 399622 256294 399678 256350
rect 399250 256170 399306 256226
rect 399374 256170 399430 256226
rect 399498 256170 399554 256226
rect 399622 256170 399678 256226
rect 399250 256046 399306 256102
rect 399374 256046 399430 256102
rect 399498 256046 399554 256102
rect 399622 256046 399678 256102
rect 399250 255922 399306 255978
rect 399374 255922 399430 255978
rect 399498 255922 399554 255978
rect 399622 255922 399678 255978
rect 384970 244294 385026 244350
rect 385094 244294 385150 244350
rect 385218 244294 385274 244350
rect 385342 244294 385398 244350
rect 384970 244170 385026 244226
rect 385094 244170 385150 244226
rect 385218 244170 385274 244226
rect 385342 244170 385398 244226
rect 384970 244046 385026 244102
rect 385094 244046 385150 244102
rect 385218 244046 385274 244102
rect 385342 244046 385398 244102
rect 384970 243922 385026 243978
rect 385094 243922 385150 243978
rect 385218 243922 385274 243978
rect 385342 243922 385398 243978
rect 387078 244294 387134 244350
rect 387202 244294 387258 244350
rect 387078 244170 387134 244226
rect 387202 244170 387258 244226
rect 387078 244046 387134 244102
rect 387202 244046 387258 244102
rect 387078 243922 387134 243978
rect 387202 243922 387258 243978
rect 402438 256294 402494 256350
rect 402562 256294 402618 256350
rect 402438 256170 402494 256226
rect 402562 256170 402618 256226
rect 402438 256046 402494 256102
rect 402562 256046 402618 256102
rect 402438 255922 402494 255978
rect 402562 255922 402618 255978
rect 417798 262294 417854 262350
rect 417922 262294 417978 262350
rect 417798 262170 417854 262226
rect 417922 262170 417978 262226
rect 417798 262046 417854 262102
rect 417922 262046 417978 262102
rect 417798 261922 417854 261978
rect 417922 261922 417978 261978
rect 433158 274294 433214 274350
rect 433282 274294 433338 274350
rect 433158 274170 433214 274226
rect 433282 274170 433338 274226
rect 433158 274046 433214 274102
rect 433282 274046 433338 274102
rect 433158 273922 433214 273978
rect 433282 273922 433338 273978
rect 435250 274294 435306 274350
rect 435374 274294 435430 274350
rect 435498 274294 435554 274350
rect 435622 274294 435678 274350
rect 435250 274170 435306 274226
rect 435374 274170 435430 274226
rect 435498 274170 435554 274226
rect 435622 274170 435678 274226
rect 435250 274046 435306 274102
rect 435374 274046 435430 274102
rect 435498 274046 435554 274102
rect 435622 274046 435678 274102
rect 435250 273922 435306 273978
rect 435374 273922 435430 273978
rect 435498 273922 435554 273978
rect 435622 273922 435678 273978
rect 420970 262294 421026 262350
rect 421094 262294 421150 262350
rect 421218 262294 421274 262350
rect 421342 262294 421398 262350
rect 420970 262170 421026 262226
rect 421094 262170 421150 262226
rect 421218 262170 421274 262226
rect 421342 262170 421398 262226
rect 420970 262046 421026 262102
rect 421094 262046 421150 262102
rect 421218 262046 421274 262102
rect 421342 262046 421398 262102
rect 420970 261922 421026 261978
rect 421094 261922 421150 261978
rect 421218 261922 421274 261978
rect 421342 261922 421398 261978
rect 402970 244294 403026 244350
rect 403094 244294 403150 244350
rect 403218 244294 403274 244350
rect 403342 244294 403398 244350
rect 402970 244170 403026 244226
rect 403094 244170 403150 244226
rect 403218 244170 403274 244226
rect 403342 244170 403398 244226
rect 402970 244046 403026 244102
rect 403094 244046 403150 244102
rect 403218 244046 403274 244102
rect 403342 244046 403398 244102
rect 402970 243922 403026 243978
rect 403094 243922 403150 243978
rect 403218 243922 403274 243978
rect 403342 243922 403398 243978
rect 399250 238294 399306 238350
rect 399374 238294 399430 238350
rect 399498 238294 399554 238350
rect 399622 238294 399678 238350
rect 399250 238170 399306 238226
rect 399374 238170 399430 238226
rect 399498 238170 399554 238226
rect 399622 238170 399678 238226
rect 399250 238046 399306 238102
rect 399374 238046 399430 238102
rect 399498 238046 399554 238102
rect 399622 238046 399678 238102
rect 399250 237922 399306 237978
rect 399374 237922 399430 237978
rect 399498 237922 399554 237978
rect 399622 237922 399678 237978
rect 384970 226294 385026 226350
rect 385094 226294 385150 226350
rect 385218 226294 385274 226350
rect 385342 226294 385398 226350
rect 384970 226170 385026 226226
rect 385094 226170 385150 226226
rect 385218 226170 385274 226226
rect 385342 226170 385398 226226
rect 384970 226046 385026 226102
rect 385094 226046 385150 226102
rect 385218 226046 385274 226102
rect 385342 226046 385398 226102
rect 384970 225922 385026 225978
rect 385094 225922 385150 225978
rect 385218 225922 385274 225978
rect 385342 225922 385398 225978
rect 387078 226294 387134 226350
rect 387202 226294 387258 226350
rect 387078 226170 387134 226226
rect 387202 226170 387258 226226
rect 387078 226046 387134 226102
rect 387202 226046 387258 226102
rect 387078 225922 387134 225978
rect 387202 225922 387258 225978
rect 402438 238294 402494 238350
rect 402562 238294 402618 238350
rect 402438 238170 402494 238226
rect 402562 238170 402618 238226
rect 402438 238046 402494 238102
rect 402562 238046 402618 238102
rect 402438 237922 402494 237978
rect 402562 237922 402618 237978
rect 417798 244294 417854 244350
rect 417922 244294 417978 244350
rect 417798 244170 417854 244226
rect 417922 244170 417978 244226
rect 417798 244046 417854 244102
rect 417922 244046 417978 244102
rect 417798 243922 417854 243978
rect 417922 243922 417978 243978
rect 433158 256294 433214 256350
rect 433282 256294 433338 256350
rect 433158 256170 433214 256226
rect 433282 256170 433338 256226
rect 433158 256046 433214 256102
rect 433282 256046 433338 256102
rect 433158 255922 433214 255978
rect 433282 255922 433338 255978
rect 435250 256294 435306 256350
rect 435374 256294 435430 256350
rect 435498 256294 435554 256350
rect 435622 256294 435678 256350
rect 435250 256170 435306 256226
rect 435374 256170 435430 256226
rect 435498 256170 435554 256226
rect 435622 256170 435678 256226
rect 435250 256046 435306 256102
rect 435374 256046 435430 256102
rect 435498 256046 435554 256102
rect 435622 256046 435678 256102
rect 435250 255922 435306 255978
rect 435374 255922 435430 255978
rect 435498 255922 435554 255978
rect 435622 255922 435678 255978
rect 420970 244294 421026 244350
rect 421094 244294 421150 244350
rect 421218 244294 421274 244350
rect 421342 244294 421398 244350
rect 420970 244170 421026 244226
rect 421094 244170 421150 244226
rect 421218 244170 421274 244226
rect 421342 244170 421398 244226
rect 420970 244046 421026 244102
rect 421094 244046 421150 244102
rect 421218 244046 421274 244102
rect 421342 244046 421398 244102
rect 420970 243922 421026 243978
rect 421094 243922 421150 243978
rect 421218 243922 421274 243978
rect 421342 243922 421398 243978
rect 402970 226294 403026 226350
rect 403094 226294 403150 226350
rect 403218 226294 403274 226350
rect 403342 226294 403398 226350
rect 402970 226170 403026 226226
rect 403094 226170 403150 226226
rect 403218 226170 403274 226226
rect 403342 226170 403398 226226
rect 402970 226046 403026 226102
rect 403094 226046 403150 226102
rect 403218 226046 403274 226102
rect 403342 226046 403398 226102
rect 402970 225922 403026 225978
rect 403094 225922 403150 225978
rect 403218 225922 403274 225978
rect 403342 225922 403398 225978
rect 399250 220294 399306 220350
rect 399374 220294 399430 220350
rect 399498 220294 399554 220350
rect 399622 220294 399678 220350
rect 399250 220170 399306 220226
rect 399374 220170 399430 220226
rect 399498 220170 399554 220226
rect 399622 220170 399678 220226
rect 399250 220046 399306 220102
rect 399374 220046 399430 220102
rect 399498 220046 399554 220102
rect 399622 220046 399678 220102
rect 399250 219922 399306 219978
rect 399374 219922 399430 219978
rect 399498 219922 399554 219978
rect 399622 219922 399678 219978
rect 384970 208294 385026 208350
rect 385094 208294 385150 208350
rect 385218 208294 385274 208350
rect 385342 208294 385398 208350
rect 384970 208170 385026 208226
rect 385094 208170 385150 208226
rect 385218 208170 385274 208226
rect 385342 208170 385398 208226
rect 384970 208046 385026 208102
rect 385094 208046 385150 208102
rect 385218 208046 385274 208102
rect 385342 208046 385398 208102
rect 384970 207922 385026 207978
rect 385094 207922 385150 207978
rect 385218 207922 385274 207978
rect 385342 207922 385398 207978
rect 387078 208294 387134 208350
rect 387202 208294 387258 208350
rect 387078 208170 387134 208226
rect 387202 208170 387258 208226
rect 387078 208046 387134 208102
rect 387202 208046 387258 208102
rect 387078 207922 387134 207978
rect 387202 207922 387258 207978
rect 402438 220294 402494 220350
rect 402562 220294 402618 220350
rect 402438 220170 402494 220226
rect 402562 220170 402618 220226
rect 402438 220046 402494 220102
rect 402562 220046 402618 220102
rect 402438 219922 402494 219978
rect 402562 219922 402618 219978
rect 417798 226294 417854 226350
rect 417922 226294 417978 226350
rect 417798 226170 417854 226226
rect 417922 226170 417978 226226
rect 417798 226046 417854 226102
rect 417922 226046 417978 226102
rect 417798 225922 417854 225978
rect 417922 225922 417978 225978
rect 433158 238294 433214 238350
rect 433282 238294 433338 238350
rect 433158 238170 433214 238226
rect 433282 238170 433338 238226
rect 433158 238046 433214 238102
rect 433282 238046 433338 238102
rect 433158 237922 433214 237978
rect 433282 237922 433338 237978
rect 435250 238294 435306 238350
rect 435374 238294 435430 238350
rect 435498 238294 435554 238350
rect 435622 238294 435678 238350
rect 435250 238170 435306 238226
rect 435374 238170 435430 238226
rect 435498 238170 435554 238226
rect 435622 238170 435678 238226
rect 435250 238046 435306 238102
rect 435374 238046 435430 238102
rect 435498 238046 435554 238102
rect 435622 238046 435678 238102
rect 435250 237922 435306 237978
rect 435374 237922 435430 237978
rect 435498 237922 435554 237978
rect 435622 237922 435678 237978
rect 420970 226294 421026 226350
rect 421094 226294 421150 226350
rect 421218 226294 421274 226350
rect 421342 226294 421398 226350
rect 420970 226170 421026 226226
rect 421094 226170 421150 226226
rect 421218 226170 421274 226226
rect 421342 226170 421398 226226
rect 420970 226046 421026 226102
rect 421094 226046 421150 226102
rect 421218 226046 421274 226102
rect 421342 226046 421398 226102
rect 420970 225922 421026 225978
rect 421094 225922 421150 225978
rect 421218 225922 421274 225978
rect 421342 225922 421398 225978
rect 402970 208294 403026 208350
rect 403094 208294 403150 208350
rect 403218 208294 403274 208350
rect 403342 208294 403398 208350
rect 402970 208170 403026 208226
rect 403094 208170 403150 208226
rect 403218 208170 403274 208226
rect 403342 208170 403398 208226
rect 402970 208046 403026 208102
rect 403094 208046 403150 208102
rect 403218 208046 403274 208102
rect 403342 208046 403398 208102
rect 402970 207922 403026 207978
rect 403094 207922 403150 207978
rect 403218 207922 403274 207978
rect 403342 207922 403398 207978
rect 399250 202294 399306 202350
rect 399374 202294 399430 202350
rect 399498 202294 399554 202350
rect 399622 202294 399678 202350
rect 399250 202170 399306 202226
rect 399374 202170 399430 202226
rect 399498 202170 399554 202226
rect 399622 202170 399678 202226
rect 399250 202046 399306 202102
rect 399374 202046 399430 202102
rect 399498 202046 399554 202102
rect 399622 202046 399678 202102
rect 399250 201922 399306 201978
rect 399374 201922 399430 201978
rect 399498 201922 399554 201978
rect 399622 201922 399678 201978
rect 384970 190294 385026 190350
rect 385094 190294 385150 190350
rect 385218 190294 385274 190350
rect 385342 190294 385398 190350
rect 384970 190170 385026 190226
rect 385094 190170 385150 190226
rect 385218 190170 385274 190226
rect 385342 190170 385398 190226
rect 384970 190046 385026 190102
rect 385094 190046 385150 190102
rect 385218 190046 385274 190102
rect 385342 190046 385398 190102
rect 384970 189922 385026 189978
rect 385094 189922 385150 189978
rect 385218 189922 385274 189978
rect 385342 189922 385398 189978
rect 387078 190294 387134 190350
rect 387202 190294 387258 190350
rect 387078 190170 387134 190226
rect 387202 190170 387258 190226
rect 387078 190046 387134 190102
rect 387202 190046 387258 190102
rect 387078 189922 387134 189978
rect 387202 189922 387258 189978
rect 402438 202294 402494 202350
rect 402562 202294 402618 202350
rect 402438 202170 402494 202226
rect 402562 202170 402618 202226
rect 402438 202046 402494 202102
rect 402562 202046 402618 202102
rect 402438 201922 402494 201978
rect 402562 201922 402618 201978
rect 417798 208294 417854 208350
rect 417922 208294 417978 208350
rect 417798 208170 417854 208226
rect 417922 208170 417978 208226
rect 417798 208046 417854 208102
rect 417922 208046 417978 208102
rect 417798 207922 417854 207978
rect 417922 207922 417978 207978
rect 433158 220294 433214 220350
rect 433282 220294 433338 220350
rect 433158 220170 433214 220226
rect 433282 220170 433338 220226
rect 433158 220046 433214 220102
rect 433282 220046 433338 220102
rect 433158 219922 433214 219978
rect 433282 219922 433338 219978
rect 435250 220294 435306 220350
rect 435374 220294 435430 220350
rect 435498 220294 435554 220350
rect 435622 220294 435678 220350
rect 435250 220170 435306 220226
rect 435374 220170 435430 220226
rect 435498 220170 435554 220226
rect 435622 220170 435678 220226
rect 435250 220046 435306 220102
rect 435374 220046 435430 220102
rect 435498 220046 435554 220102
rect 435622 220046 435678 220102
rect 435250 219922 435306 219978
rect 435374 219922 435430 219978
rect 435498 219922 435554 219978
rect 435622 219922 435678 219978
rect 420970 208294 421026 208350
rect 421094 208294 421150 208350
rect 421218 208294 421274 208350
rect 421342 208294 421398 208350
rect 420970 208170 421026 208226
rect 421094 208170 421150 208226
rect 421218 208170 421274 208226
rect 421342 208170 421398 208226
rect 420970 208046 421026 208102
rect 421094 208046 421150 208102
rect 421218 208046 421274 208102
rect 421342 208046 421398 208102
rect 420970 207922 421026 207978
rect 421094 207922 421150 207978
rect 421218 207922 421274 207978
rect 421342 207922 421398 207978
rect 402970 190294 403026 190350
rect 403094 190294 403150 190350
rect 403218 190294 403274 190350
rect 403342 190294 403398 190350
rect 402970 190170 403026 190226
rect 403094 190170 403150 190226
rect 403218 190170 403274 190226
rect 403342 190170 403398 190226
rect 402970 190046 403026 190102
rect 403094 190046 403150 190102
rect 403218 190046 403274 190102
rect 403342 190046 403398 190102
rect 402970 189922 403026 189978
rect 403094 189922 403150 189978
rect 403218 189922 403274 189978
rect 403342 189922 403398 189978
rect 399250 184294 399306 184350
rect 399374 184294 399430 184350
rect 399498 184294 399554 184350
rect 399622 184294 399678 184350
rect 399250 184170 399306 184226
rect 399374 184170 399430 184226
rect 399498 184170 399554 184226
rect 399622 184170 399678 184226
rect 399250 184046 399306 184102
rect 399374 184046 399430 184102
rect 399498 184046 399554 184102
rect 399622 184046 399678 184102
rect 399250 183922 399306 183978
rect 399374 183922 399430 183978
rect 399498 183922 399554 183978
rect 399622 183922 399678 183978
rect 384970 172294 385026 172350
rect 385094 172294 385150 172350
rect 385218 172294 385274 172350
rect 385342 172294 385398 172350
rect 384970 172170 385026 172226
rect 385094 172170 385150 172226
rect 385218 172170 385274 172226
rect 385342 172170 385398 172226
rect 384970 172046 385026 172102
rect 385094 172046 385150 172102
rect 385218 172046 385274 172102
rect 385342 172046 385398 172102
rect 384970 171922 385026 171978
rect 385094 171922 385150 171978
rect 385218 171922 385274 171978
rect 385342 171922 385398 171978
rect 387078 172294 387134 172350
rect 387202 172294 387258 172350
rect 387078 172170 387134 172226
rect 387202 172170 387258 172226
rect 387078 172046 387134 172102
rect 387202 172046 387258 172102
rect 387078 171922 387134 171978
rect 387202 171922 387258 171978
rect 402438 184294 402494 184350
rect 402562 184294 402618 184350
rect 402438 184170 402494 184226
rect 402562 184170 402618 184226
rect 402438 184046 402494 184102
rect 402562 184046 402618 184102
rect 402438 183922 402494 183978
rect 402562 183922 402618 183978
rect 417798 190294 417854 190350
rect 417922 190294 417978 190350
rect 417798 190170 417854 190226
rect 417922 190170 417978 190226
rect 417798 190046 417854 190102
rect 417922 190046 417978 190102
rect 417798 189922 417854 189978
rect 417922 189922 417978 189978
rect 433158 202294 433214 202350
rect 433282 202294 433338 202350
rect 433158 202170 433214 202226
rect 433282 202170 433338 202226
rect 433158 202046 433214 202102
rect 433282 202046 433338 202102
rect 433158 201922 433214 201978
rect 433282 201922 433338 201978
rect 435250 202294 435306 202350
rect 435374 202294 435430 202350
rect 435498 202294 435554 202350
rect 435622 202294 435678 202350
rect 435250 202170 435306 202226
rect 435374 202170 435430 202226
rect 435498 202170 435554 202226
rect 435622 202170 435678 202226
rect 435250 202046 435306 202102
rect 435374 202046 435430 202102
rect 435498 202046 435554 202102
rect 435622 202046 435678 202102
rect 435250 201922 435306 201978
rect 435374 201922 435430 201978
rect 435498 201922 435554 201978
rect 435622 201922 435678 201978
rect 420970 190294 421026 190350
rect 421094 190294 421150 190350
rect 421218 190294 421274 190350
rect 421342 190294 421398 190350
rect 420970 190170 421026 190226
rect 421094 190170 421150 190226
rect 421218 190170 421274 190226
rect 421342 190170 421398 190226
rect 420970 190046 421026 190102
rect 421094 190046 421150 190102
rect 421218 190046 421274 190102
rect 421342 190046 421398 190102
rect 420970 189922 421026 189978
rect 421094 189922 421150 189978
rect 421218 189922 421274 189978
rect 421342 189922 421398 189978
rect 402970 172294 403026 172350
rect 403094 172294 403150 172350
rect 403218 172294 403274 172350
rect 403342 172294 403398 172350
rect 402970 172170 403026 172226
rect 403094 172170 403150 172226
rect 403218 172170 403274 172226
rect 403342 172170 403398 172226
rect 402970 172046 403026 172102
rect 403094 172046 403150 172102
rect 403218 172046 403274 172102
rect 403342 172046 403398 172102
rect 402970 171922 403026 171978
rect 403094 171922 403150 171978
rect 403218 171922 403274 171978
rect 403342 171922 403398 171978
rect 399250 166294 399306 166350
rect 399374 166294 399430 166350
rect 399498 166294 399554 166350
rect 399622 166294 399678 166350
rect 399250 166170 399306 166226
rect 399374 166170 399430 166226
rect 399498 166170 399554 166226
rect 399622 166170 399678 166226
rect 399250 166046 399306 166102
rect 399374 166046 399430 166102
rect 399498 166046 399554 166102
rect 399622 166046 399678 166102
rect 399250 165922 399306 165978
rect 399374 165922 399430 165978
rect 399498 165922 399554 165978
rect 399622 165922 399678 165978
rect 384970 154294 385026 154350
rect 385094 154294 385150 154350
rect 385218 154294 385274 154350
rect 385342 154294 385398 154350
rect 384970 154170 385026 154226
rect 385094 154170 385150 154226
rect 385218 154170 385274 154226
rect 385342 154170 385398 154226
rect 384970 154046 385026 154102
rect 385094 154046 385150 154102
rect 385218 154046 385274 154102
rect 385342 154046 385398 154102
rect 384970 153922 385026 153978
rect 385094 153922 385150 153978
rect 385218 153922 385274 153978
rect 385342 153922 385398 153978
rect 387078 154294 387134 154350
rect 387202 154294 387258 154350
rect 387078 154170 387134 154226
rect 387202 154170 387258 154226
rect 387078 154046 387134 154102
rect 387202 154046 387258 154102
rect 387078 153922 387134 153978
rect 387202 153922 387258 153978
rect 402438 166294 402494 166350
rect 402562 166294 402618 166350
rect 402438 166170 402494 166226
rect 402562 166170 402618 166226
rect 402438 166046 402494 166102
rect 402562 166046 402618 166102
rect 402438 165922 402494 165978
rect 402562 165922 402618 165978
rect 417798 172294 417854 172350
rect 417922 172294 417978 172350
rect 417798 172170 417854 172226
rect 417922 172170 417978 172226
rect 417798 172046 417854 172102
rect 417922 172046 417978 172102
rect 417798 171922 417854 171978
rect 417922 171922 417978 171978
rect 433158 184294 433214 184350
rect 433282 184294 433338 184350
rect 433158 184170 433214 184226
rect 433282 184170 433338 184226
rect 433158 184046 433214 184102
rect 433282 184046 433338 184102
rect 433158 183922 433214 183978
rect 433282 183922 433338 183978
rect 435250 184294 435306 184350
rect 435374 184294 435430 184350
rect 435498 184294 435554 184350
rect 435622 184294 435678 184350
rect 435250 184170 435306 184226
rect 435374 184170 435430 184226
rect 435498 184170 435554 184226
rect 435622 184170 435678 184226
rect 435250 184046 435306 184102
rect 435374 184046 435430 184102
rect 435498 184046 435554 184102
rect 435622 184046 435678 184102
rect 435250 183922 435306 183978
rect 435374 183922 435430 183978
rect 435498 183922 435554 183978
rect 435622 183922 435678 183978
rect 420970 172294 421026 172350
rect 421094 172294 421150 172350
rect 421218 172294 421274 172350
rect 421342 172294 421398 172350
rect 420970 172170 421026 172226
rect 421094 172170 421150 172226
rect 421218 172170 421274 172226
rect 421342 172170 421398 172226
rect 420970 172046 421026 172102
rect 421094 172046 421150 172102
rect 421218 172046 421274 172102
rect 421342 172046 421398 172102
rect 420970 171922 421026 171978
rect 421094 171922 421150 171978
rect 421218 171922 421274 171978
rect 421342 171922 421398 171978
rect 402970 154294 403026 154350
rect 403094 154294 403150 154350
rect 403218 154294 403274 154350
rect 403342 154294 403398 154350
rect 402970 154170 403026 154226
rect 403094 154170 403150 154226
rect 403218 154170 403274 154226
rect 403342 154170 403398 154226
rect 402970 154046 403026 154102
rect 403094 154046 403150 154102
rect 403218 154046 403274 154102
rect 403342 154046 403398 154102
rect 402970 153922 403026 153978
rect 403094 153922 403150 153978
rect 403218 153922 403274 153978
rect 403342 153922 403398 153978
rect 399250 148294 399306 148350
rect 399374 148294 399430 148350
rect 399498 148294 399554 148350
rect 399622 148294 399678 148350
rect 399250 148170 399306 148226
rect 399374 148170 399430 148226
rect 399498 148170 399554 148226
rect 399622 148170 399678 148226
rect 399250 148046 399306 148102
rect 399374 148046 399430 148102
rect 399498 148046 399554 148102
rect 399622 148046 399678 148102
rect 399250 147922 399306 147978
rect 399374 147922 399430 147978
rect 399498 147922 399554 147978
rect 399622 147922 399678 147978
rect 384970 136294 385026 136350
rect 385094 136294 385150 136350
rect 385218 136294 385274 136350
rect 385342 136294 385398 136350
rect 384970 136170 385026 136226
rect 385094 136170 385150 136226
rect 385218 136170 385274 136226
rect 385342 136170 385398 136226
rect 384970 136046 385026 136102
rect 385094 136046 385150 136102
rect 385218 136046 385274 136102
rect 385342 136046 385398 136102
rect 384970 135922 385026 135978
rect 385094 135922 385150 135978
rect 385218 135922 385274 135978
rect 385342 135922 385398 135978
rect 387078 136294 387134 136350
rect 387202 136294 387258 136350
rect 387078 136170 387134 136226
rect 387202 136170 387258 136226
rect 387078 136046 387134 136102
rect 387202 136046 387258 136102
rect 387078 135922 387134 135978
rect 387202 135922 387258 135978
rect 402438 148294 402494 148350
rect 402562 148294 402618 148350
rect 402438 148170 402494 148226
rect 402562 148170 402618 148226
rect 402438 148046 402494 148102
rect 402562 148046 402618 148102
rect 402438 147922 402494 147978
rect 402562 147922 402618 147978
rect 417798 154294 417854 154350
rect 417922 154294 417978 154350
rect 417798 154170 417854 154226
rect 417922 154170 417978 154226
rect 417798 154046 417854 154102
rect 417922 154046 417978 154102
rect 417798 153922 417854 153978
rect 417922 153922 417978 153978
rect 433158 166294 433214 166350
rect 433282 166294 433338 166350
rect 433158 166170 433214 166226
rect 433282 166170 433338 166226
rect 433158 166046 433214 166102
rect 433282 166046 433338 166102
rect 433158 165922 433214 165978
rect 433282 165922 433338 165978
rect 435250 166294 435306 166350
rect 435374 166294 435430 166350
rect 435498 166294 435554 166350
rect 435622 166294 435678 166350
rect 435250 166170 435306 166226
rect 435374 166170 435430 166226
rect 435498 166170 435554 166226
rect 435622 166170 435678 166226
rect 435250 166046 435306 166102
rect 435374 166046 435430 166102
rect 435498 166046 435554 166102
rect 435622 166046 435678 166102
rect 435250 165922 435306 165978
rect 435374 165922 435430 165978
rect 435498 165922 435554 165978
rect 435622 165922 435678 165978
rect 420970 154294 421026 154350
rect 421094 154294 421150 154350
rect 421218 154294 421274 154350
rect 421342 154294 421398 154350
rect 420970 154170 421026 154226
rect 421094 154170 421150 154226
rect 421218 154170 421274 154226
rect 421342 154170 421398 154226
rect 420970 154046 421026 154102
rect 421094 154046 421150 154102
rect 421218 154046 421274 154102
rect 421342 154046 421398 154102
rect 420970 153922 421026 153978
rect 421094 153922 421150 153978
rect 421218 153922 421274 153978
rect 421342 153922 421398 153978
rect 402970 136294 403026 136350
rect 403094 136294 403150 136350
rect 403218 136294 403274 136350
rect 403342 136294 403398 136350
rect 402970 136170 403026 136226
rect 403094 136170 403150 136226
rect 403218 136170 403274 136226
rect 403342 136170 403398 136226
rect 402970 136046 403026 136102
rect 403094 136046 403150 136102
rect 403218 136046 403274 136102
rect 403342 136046 403398 136102
rect 402970 135922 403026 135978
rect 403094 135922 403150 135978
rect 403218 135922 403274 135978
rect 403342 135922 403398 135978
rect 399250 130294 399306 130350
rect 399374 130294 399430 130350
rect 399498 130294 399554 130350
rect 399622 130294 399678 130350
rect 399250 130170 399306 130226
rect 399374 130170 399430 130226
rect 399498 130170 399554 130226
rect 399622 130170 399678 130226
rect 399250 130046 399306 130102
rect 399374 130046 399430 130102
rect 399498 130046 399554 130102
rect 399622 130046 399678 130102
rect 399250 129922 399306 129978
rect 399374 129922 399430 129978
rect 399498 129922 399554 129978
rect 399622 129922 399678 129978
rect 384970 118294 385026 118350
rect 385094 118294 385150 118350
rect 385218 118294 385274 118350
rect 385342 118294 385398 118350
rect 384970 118170 385026 118226
rect 385094 118170 385150 118226
rect 385218 118170 385274 118226
rect 385342 118170 385398 118226
rect 384970 118046 385026 118102
rect 385094 118046 385150 118102
rect 385218 118046 385274 118102
rect 385342 118046 385398 118102
rect 384970 117922 385026 117978
rect 385094 117922 385150 117978
rect 385218 117922 385274 117978
rect 385342 117922 385398 117978
rect 387078 118294 387134 118350
rect 387202 118294 387258 118350
rect 387078 118170 387134 118226
rect 387202 118170 387258 118226
rect 387078 118046 387134 118102
rect 387202 118046 387258 118102
rect 387078 117922 387134 117978
rect 387202 117922 387258 117978
rect 402438 130294 402494 130350
rect 402562 130294 402618 130350
rect 402438 130170 402494 130226
rect 402562 130170 402618 130226
rect 402438 130046 402494 130102
rect 402562 130046 402618 130102
rect 402438 129922 402494 129978
rect 402562 129922 402618 129978
rect 417798 136294 417854 136350
rect 417922 136294 417978 136350
rect 417798 136170 417854 136226
rect 417922 136170 417978 136226
rect 417798 136046 417854 136102
rect 417922 136046 417978 136102
rect 417798 135922 417854 135978
rect 417922 135922 417978 135978
rect 433158 148294 433214 148350
rect 433282 148294 433338 148350
rect 433158 148170 433214 148226
rect 433282 148170 433338 148226
rect 433158 148046 433214 148102
rect 433282 148046 433338 148102
rect 433158 147922 433214 147978
rect 433282 147922 433338 147978
rect 435250 148294 435306 148350
rect 435374 148294 435430 148350
rect 435498 148294 435554 148350
rect 435622 148294 435678 148350
rect 435250 148170 435306 148226
rect 435374 148170 435430 148226
rect 435498 148170 435554 148226
rect 435622 148170 435678 148226
rect 435250 148046 435306 148102
rect 435374 148046 435430 148102
rect 435498 148046 435554 148102
rect 435622 148046 435678 148102
rect 435250 147922 435306 147978
rect 435374 147922 435430 147978
rect 435498 147922 435554 147978
rect 435622 147922 435678 147978
rect 420970 136294 421026 136350
rect 421094 136294 421150 136350
rect 421218 136294 421274 136350
rect 421342 136294 421398 136350
rect 420970 136170 421026 136226
rect 421094 136170 421150 136226
rect 421218 136170 421274 136226
rect 421342 136170 421398 136226
rect 420970 136046 421026 136102
rect 421094 136046 421150 136102
rect 421218 136046 421274 136102
rect 421342 136046 421398 136102
rect 420970 135922 421026 135978
rect 421094 135922 421150 135978
rect 421218 135922 421274 135978
rect 421342 135922 421398 135978
rect 402970 118294 403026 118350
rect 403094 118294 403150 118350
rect 403218 118294 403274 118350
rect 403342 118294 403398 118350
rect 402970 118170 403026 118226
rect 403094 118170 403150 118226
rect 403218 118170 403274 118226
rect 403342 118170 403398 118226
rect 402970 118046 403026 118102
rect 403094 118046 403150 118102
rect 403218 118046 403274 118102
rect 403342 118046 403398 118102
rect 402970 117922 403026 117978
rect 403094 117922 403150 117978
rect 403218 117922 403274 117978
rect 403342 117922 403398 117978
rect 399250 112294 399306 112350
rect 399374 112294 399430 112350
rect 399498 112294 399554 112350
rect 399622 112294 399678 112350
rect 399250 112170 399306 112226
rect 399374 112170 399430 112226
rect 399498 112170 399554 112226
rect 399622 112170 399678 112226
rect 399250 112046 399306 112102
rect 399374 112046 399430 112102
rect 399498 112046 399554 112102
rect 399622 112046 399678 112102
rect 399250 111922 399306 111978
rect 399374 111922 399430 111978
rect 399498 111922 399554 111978
rect 399622 111922 399678 111978
rect 384970 100294 385026 100350
rect 385094 100294 385150 100350
rect 385218 100294 385274 100350
rect 385342 100294 385398 100350
rect 384970 100170 385026 100226
rect 385094 100170 385150 100226
rect 385218 100170 385274 100226
rect 385342 100170 385398 100226
rect 384970 100046 385026 100102
rect 385094 100046 385150 100102
rect 385218 100046 385274 100102
rect 385342 100046 385398 100102
rect 384970 99922 385026 99978
rect 385094 99922 385150 99978
rect 385218 99922 385274 99978
rect 385342 99922 385398 99978
rect 387078 100294 387134 100350
rect 387202 100294 387258 100350
rect 387078 100170 387134 100226
rect 387202 100170 387258 100226
rect 387078 100046 387134 100102
rect 387202 100046 387258 100102
rect 387078 99922 387134 99978
rect 387202 99922 387258 99978
rect 402438 112294 402494 112350
rect 402562 112294 402618 112350
rect 402438 112170 402494 112226
rect 402562 112170 402618 112226
rect 402438 112046 402494 112102
rect 402562 112046 402618 112102
rect 402438 111922 402494 111978
rect 402562 111922 402618 111978
rect 417798 118294 417854 118350
rect 417922 118294 417978 118350
rect 417798 118170 417854 118226
rect 417922 118170 417978 118226
rect 417798 118046 417854 118102
rect 417922 118046 417978 118102
rect 417798 117922 417854 117978
rect 417922 117922 417978 117978
rect 433158 130294 433214 130350
rect 433282 130294 433338 130350
rect 433158 130170 433214 130226
rect 433282 130170 433338 130226
rect 433158 130046 433214 130102
rect 433282 130046 433338 130102
rect 433158 129922 433214 129978
rect 433282 129922 433338 129978
rect 435250 130294 435306 130350
rect 435374 130294 435430 130350
rect 435498 130294 435554 130350
rect 435622 130294 435678 130350
rect 435250 130170 435306 130226
rect 435374 130170 435430 130226
rect 435498 130170 435554 130226
rect 435622 130170 435678 130226
rect 435250 130046 435306 130102
rect 435374 130046 435430 130102
rect 435498 130046 435554 130102
rect 435622 130046 435678 130102
rect 435250 129922 435306 129978
rect 435374 129922 435430 129978
rect 435498 129922 435554 129978
rect 435622 129922 435678 129978
rect 420970 118294 421026 118350
rect 421094 118294 421150 118350
rect 421218 118294 421274 118350
rect 421342 118294 421398 118350
rect 420970 118170 421026 118226
rect 421094 118170 421150 118226
rect 421218 118170 421274 118226
rect 421342 118170 421398 118226
rect 420970 118046 421026 118102
rect 421094 118046 421150 118102
rect 421218 118046 421274 118102
rect 421342 118046 421398 118102
rect 420970 117922 421026 117978
rect 421094 117922 421150 117978
rect 421218 117922 421274 117978
rect 421342 117922 421398 117978
rect 402970 100294 403026 100350
rect 403094 100294 403150 100350
rect 403218 100294 403274 100350
rect 403342 100294 403398 100350
rect 402970 100170 403026 100226
rect 403094 100170 403150 100226
rect 403218 100170 403274 100226
rect 403342 100170 403398 100226
rect 402970 100046 403026 100102
rect 403094 100046 403150 100102
rect 403218 100046 403274 100102
rect 403342 100046 403398 100102
rect 402970 99922 403026 99978
rect 403094 99922 403150 99978
rect 403218 99922 403274 99978
rect 403342 99922 403398 99978
rect 399250 94294 399306 94350
rect 399374 94294 399430 94350
rect 399498 94294 399554 94350
rect 399622 94294 399678 94350
rect 399250 94170 399306 94226
rect 399374 94170 399430 94226
rect 399498 94170 399554 94226
rect 399622 94170 399678 94226
rect 399250 94046 399306 94102
rect 399374 94046 399430 94102
rect 399498 94046 399554 94102
rect 399622 94046 399678 94102
rect 399250 93922 399306 93978
rect 399374 93922 399430 93978
rect 399498 93922 399554 93978
rect 399622 93922 399678 93978
rect 384970 82294 385026 82350
rect 385094 82294 385150 82350
rect 385218 82294 385274 82350
rect 385342 82294 385398 82350
rect 384970 82170 385026 82226
rect 385094 82170 385150 82226
rect 385218 82170 385274 82226
rect 385342 82170 385398 82226
rect 384970 82046 385026 82102
rect 385094 82046 385150 82102
rect 385218 82046 385274 82102
rect 385342 82046 385398 82102
rect 384970 81922 385026 81978
rect 385094 81922 385150 81978
rect 385218 81922 385274 81978
rect 385342 81922 385398 81978
rect 387078 82294 387134 82350
rect 387202 82294 387258 82350
rect 387078 82170 387134 82226
rect 387202 82170 387258 82226
rect 387078 82046 387134 82102
rect 387202 82046 387258 82102
rect 387078 81922 387134 81978
rect 387202 81922 387258 81978
rect 402438 94294 402494 94350
rect 402562 94294 402618 94350
rect 402438 94170 402494 94226
rect 402562 94170 402618 94226
rect 402438 94046 402494 94102
rect 402562 94046 402618 94102
rect 402438 93922 402494 93978
rect 402562 93922 402618 93978
rect 417798 100294 417854 100350
rect 417922 100294 417978 100350
rect 417798 100170 417854 100226
rect 417922 100170 417978 100226
rect 417798 100046 417854 100102
rect 417922 100046 417978 100102
rect 417798 99922 417854 99978
rect 417922 99922 417978 99978
rect 433158 112294 433214 112350
rect 433282 112294 433338 112350
rect 433158 112170 433214 112226
rect 433282 112170 433338 112226
rect 433158 112046 433214 112102
rect 433282 112046 433338 112102
rect 433158 111922 433214 111978
rect 433282 111922 433338 111978
rect 435250 112294 435306 112350
rect 435374 112294 435430 112350
rect 435498 112294 435554 112350
rect 435622 112294 435678 112350
rect 435250 112170 435306 112226
rect 435374 112170 435430 112226
rect 435498 112170 435554 112226
rect 435622 112170 435678 112226
rect 435250 112046 435306 112102
rect 435374 112046 435430 112102
rect 435498 112046 435554 112102
rect 435622 112046 435678 112102
rect 435250 111922 435306 111978
rect 435374 111922 435430 111978
rect 435498 111922 435554 111978
rect 435622 111922 435678 111978
rect 420970 100294 421026 100350
rect 421094 100294 421150 100350
rect 421218 100294 421274 100350
rect 421342 100294 421398 100350
rect 420970 100170 421026 100226
rect 421094 100170 421150 100226
rect 421218 100170 421274 100226
rect 421342 100170 421398 100226
rect 420970 100046 421026 100102
rect 421094 100046 421150 100102
rect 421218 100046 421274 100102
rect 421342 100046 421398 100102
rect 420970 99922 421026 99978
rect 421094 99922 421150 99978
rect 421218 99922 421274 99978
rect 421342 99922 421398 99978
rect 402970 82294 403026 82350
rect 403094 82294 403150 82350
rect 403218 82294 403274 82350
rect 403342 82294 403398 82350
rect 402970 82170 403026 82226
rect 403094 82170 403150 82226
rect 403218 82170 403274 82226
rect 403342 82170 403398 82226
rect 402970 82046 403026 82102
rect 403094 82046 403150 82102
rect 403218 82046 403274 82102
rect 403342 82046 403398 82102
rect 402970 81922 403026 81978
rect 403094 81922 403150 81978
rect 403218 81922 403274 81978
rect 403342 81922 403398 81978
rect 399250 76294 399306 76350
rect 399374 76294 399430 76350
rect 399498 76294 399554 76350
rect 399622 76294 399678 76350
rect 399250 76170 399306 76226
rect 399374 76170 399430 76226
rect 399498 76170 399554 76226
rect 399622 76170 399678 76226
rect 399250 76046 399306 76102
rect 399374 76046 399430 76102
rect 399498 76046 399554 76102
rect 399622 76046 399678 76102
rect 399250 75922 399306 75978
rect 399374 75922 399430 75978
rect 399498 75922 399554 75978
rect 399622 75922 399678 75978
rect 384970 64294 385026 64350
rect 385094 64294 385150 64350
rect 385218 64294 385274 64350
rect 385342 64294 385398 64350
rect 384970 64170 385026 64226
rect 385094 64170 385150 64226
rect 385218 64170 385274 64226
rect 385342 64170 385398 64226
rect 384970 64046 385026 64102
rect 385094 64046 385150 64102
rect 385218 64046 385274 64102
rect 385342 64046 385398 64102
rect 384970 63922 385026 63978
rect 385094 63922 385150 63978
rect 385218 63922 385274 63978
rect 385342 63922 385398 63978
rect 387078 64294 387134 64350
rect 387202 64294 387258 64350
rect 387078 64170 387134 64226
rect 387202 64170 387258 64226
rect 387078 64046 387134 64102
rect 387202 64046 387258 64102
rect 387078 63922 387134 63978
rect 387202 63922 387258 63978
rect 384970 46294 385026 46350
rect 385094 46294 385150 46350
rect 385218 46294 385274 46350
rect 385342 46294 385398 46350
rect 384970 46170 385026 46226
rect 385094 46170 385150 46226
rect 385218 46170 385274 46226
rect 385342 46170 385398 46226
rect 384970 46046 385026 46102
rect 385094 46046 385150 46102
rect 385218 46046 385274 46102
rect 385342 46046 385398 46102
rect 384970 45922 385026 45978
rect 385094 45922 385150 45978
rect 385218 45922 385274 45978
rect 385342 45922 385398 45978
rect 384970 28294 385026 28350
rect 385094 28294 385150 28350
rect 385218 28294 385274 28350
rect 385342 28294 385398 28350
rect 384970 28170 385026 28226
rect 385094 28170 385150 28226
rect 385218 28170 385274 28226
rect 385342 28170 385398 28226
rect 384970 28046 385026 28102
rect 385094 28046 385150 28102
rect 385218 28046 385274 28102
rect 385342 28046 385398 28102
rect 384970 27922 385026 27978
rect 385094 27922 385150 27978
rect 385218 27922 385274 27978
rect 385342 27922 385398 27978
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 402438 76294 402494 76350
rect 402562 76294 402618 76350
rect 402438 76170 402494 76226
rect 402562 76170 402618 76226
rect 402438 76046 402494 76102
rect 402562 76046 402618 76102
rect 402438 75922 402494 75978
rect 402562 75922 402618 75978
rect 399250 58294 399306 58350
rect 399374 58294 399430 58350
rect 399498 58294 399554 58350
rect 399622 58294 399678 58350
rect 399250 58170 399306 58226
rect 399374 58170 399430 58226
rect 399498 58170 399554 58226
rect 399622 58170 399678 58226
rect 399250 58046 399306 58102
rect 399374 58046 399430 58102
rect 399498 58046 399554 58102
rect 399622 58046 399678 58102
rect 399250 57922 399306 57978
rect 399374 57922 399430 57978
rect 399498 57922 399554 57978
rect 399622 57922 399678 57978
rect 399250 40294 399306 40350
rect 399374 40294 399430 40350
rect 399498 40294 399554 40350
rect 399622 40294 399678 40350
rect 399250 40170 399306 40226
rect 399374 40170 399430 40226
rect 399498 40170 399554 40226
rect 399622 40170 399678 40226
rect 399250 40046 399306 40102
rect 399374 40046 399430 40102
rect 399498 40046 399554 40102
rect 399622 40046 399678 40102
rect 399250 39922 399306 39978
rect 399374 39922 399430 39978
rect 399498 39922 399554 39978
rect 399622 39922 399678 39978
rect 399250 22294 399306 22350
rect 399374 22294 399430 22350
rect 399498 22294 399554 22350
rect 399622 22294 399678 22350
rect 399250 22170 399306 22226
rect 399374 22170 399430 22226
rect 399498 22170 399554 22226
rect 399622 22170 399678 22226
rect 399250 22046 399306 22102
rect 399374 22046 399430 22102
rect 399498 22046 399554 22102
rect 399622 22046 399678 22102
rect 399250 21922 399306 21978
rect 399374 21922 399430 21978
rect 399498 21922 399554 21978
rect 399622 21922 399678 21978
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 417798 82294 417854 82350
rect 417922 82294 417978 82350
rect 417798 82170 417854 82226
rect 417922 82170 417978 82226
rect 417798 82046 417854 82102
rect 417922 82046 417978 82102
rect 417798 81922 417854 81978
rect 417922 81922 417978 81978
rect 433158 94294 433214 94350
rect 433282 94294 433338 94350
rect 433158 94170 433214 94226
rect 433282 94170 433338 94226
rect 433158 94046 433214 94102
rect 433282 94046 433338 94102
rect 433158 93922 433214 93978
rect 433282 93922 433338 93978
rect 435250 94294 435306 94350
rect 435374 94294 435430 94350
rect 435498 94294 435554 94350
rect 435622 94294 435678 94350
rect 435250 94170 435306 94226
rect 435374 94170 435430 94226
rect 435498 94170 435554 94226
rect 435622 94170 435678 94226
rect 435250 94046 435306 94102
rect 435374 94046 435430 94102
rect 435498 94046 435554 94102
rect 435622 94046 435678 94102
rect 435250 93922 435306 93978
rect 435374 93922 435430 93978
rect 435498 93922 435554 93978
rect 435622 93922 435678 93978
rect 420970 82294 421026 82350
rect 421094 82294 421150 82350
rect 421218 82294 421274 82350
rect 421342 82294 421398 82350
rect 420970 82170 421026 82226
rect 421094 82170 421150 82226
rect 421218 82170 421274 82226
rect 421342 82170 421398 82226
rect 420970 82046 421026 82102
rect 421094 82046 421150 82102
rect 421218 82046 421274 82102
rect 421342 82046 421398 82102
rect 420970 81922 421026 81978
rect 421094 81922 421150 81978
rect 421218 81922 421274 81978
rect 421342 81922 421398 81978
rect 402970 64294 403026 64350
rect 403094 64294 403150 64350
rect 403218 64294 403274 64350
rect 403342 64294 403398 64350
rect 402970 64170 403026 64226
rect 403094 64170 403150 64226
rect 403218 64170 403274 64226
rect 403342 64170 403398 64226
rect 402970 64046 403026 64102
rect 403094 64046 403150 64102
rect 403218 64046 403274 64102
rect 403342 64046 403398 64102
rect 402970 63922 403026 63978
rect 403094 63922 403150 63978
rect 403218 63922 403274 63978
rect 403342 63922 403398 63978
rect 417798 64294 417854 64350
rect 417922 64294 417978 64350
rect 417798 64170 417854 64226
rect 417922 64170 417978 64226
rect 417798 64046 417854 64102
rect 417922 64046 417978 64102
rect 417798 63922 417854 63978
rect 417922 63922 417978 63978
rect 433158 76294 433214 76350
rect 433282 76294 433338 76350
rect 433158 76170 433214 76226
rect 433282 76170 433338 76226
rect 433158 76046 433214 76102
rect 433282 76046 433338 76102
rect 433158 75922 433214 75978
rect 433282 75922 433338 75978
rect 435250 76294 435306 76350
rect 435374 76294 435430 76350
rect 435498 76294 435554 76350
rect 435622 76294 435678 76350
rect 435250 76170 435306 76226
rect 435374 76170 435430 76226
rect 435498 76170 435554 76226
rect 435622 76170 435678 76226
rect 435250 76046 435306 76102
rect 435374 76046 435430 76102
rect 435498 76046 435554 76102
rect 435622 76046 435678 76102
rect 435250 75922 435306 75978
rect 435374 75922 435430 75978
rect 435498 75922 435554 75978
rect 435622 75922 435678 75978
rect 420970 64294 421026 64350
rect 421094 64294 421150 64350
rect 421218 64294 421274 64350
rect 421342 64294 421398 64350
rect 420970 64170 421026 64226
rect 421094 64170 421150 64226
rect 421218 64170 421274 64226
rect 421342 64170 421398 64226
rect 420970 64046 421026 64102
rect 421094 64046 421150 64102
rect 421218 64046 421274 64102
rect 421342 64046 421398 64102
rect 420970 63922 421026 63978
rect 421094 63922 421150 63978
rect 421218 63922 421274 63978
rect 421342 63922 421398 63978
rect 402970 46294 403026 46350
rect 403094 46294 403150 46350
rect 403218 46294 403274 46350
rect 403342 46294 403398 46350
rect 402970 46170 403026 46226
rect 403094 46170 403150 46226
rect 403218 46170 403274 46226
rect 403342 46170 403398 46226
rect 402970 46046 403026 46102
rect 403094 46046 403150 46102
rect 403218 46046 403274 46102
rect 403342 46046 403398 46102
rect 402970 45922 403026 45978
rect 403094 45922 403150 45978
rect 403218 45922 403274 45978
rect 403342 45922 403398 45978
rect 402970 28294 403026 28350
rect 403094 28294 403150 28350
rect 403218 28294 403274 28350
rect 403342 28294 403398 28350
rect 402970 28170 403026 28226
rect 403094 28170 403150 28226
rect 403218 28170 403274 28226
rect 403342 28170 403398 28226
rect 402970 28046 403026 28102
rect 403094 28046 403150 28102
rect 403218 28046 403274 28102
rect 403342 28046 403398 28102
rect 402970 27922 403026 27978
rect 403094 27922 403150 27978
rect 403218 27922 403274 27978
rect 403342 27922 403398 27978
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 58294 417306 58350
rect 417374 58294 417430 58350
rect 417498 58294 417554 58350
rect 417622 58294 417678 58350
rect 417250 58170 417306 58226
rect 417374 58170 417430 58226
rect 417498 58170 417554 58226
rect 417622 58170 417678 58226
rect 417250 58046 417306 58102
rect 417374 58046 417430 58102
rect 417498 58046 417554 58102
rect 417622 58046 417678 58102
rect 417250 57922 417306 57978
rect 417374 57922 417430 57978
rect 417498 57922 417554 57978
rect 417622 57922 417678 57978
rect 417250 40294 417306 40350
rect 417374 40294 417430 40350
rect 417498 40294 417554 40350
rect 417622 40294 417678 40350
rect 417250 40170 417306 40226
rect 417374 40170 417430 40226
rect 417498 40170 417554 40226
rect 417622 40170 417678 40226
rect 417250 40046 417306 40102
rect 417374 40046 417430 40102
rect 417498 40046 417554 40102
rect 417622 40046 417678 40102
rect 417250 39922 417306 39978
rect 417374 39922 417430 39978
rect 417498 39922 417554 39978
rect 417622 39922 417678 39978
rect 417250 22294 417306 22350
rect 417374 22294 417430 22350
rect 417498 22294 417554 22350
rect 417622 22294 417678 22350
rect 417250 22170 417306 22226
rect 417374 22170 417430 22226
rect 417498 22170 417554 22226
rect 417622 22170 417678 22226
rect 417250 22046 417306 22102
rect 417374 22046 417430 22102
rect 417498 22046 417554 22102
rect 417622 22046 417678 22102
rect 417250 21922 417306 21978
rect 417374 21922 417430 21978
rect 417498 21922 417554 21978
rect 417622 21922 417678 21978
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 420970 46294 421026 46350
rect 421094 46294 421150 46350
rect 421218 46294 421274 46350
rect 421342 46294 421398 46350
rect 420970 46170 421026 46226
rect 421094 46170 421150 46226
rect 421218 46170 421274 46226
rect 421342 46170 421398 46226
rect 420970 46046 421026 46102
rect 421094 46046 421150 46102
rect 421218 46046 421274 46102
rect 421342 46046 421398 46102
rect 420970 45922 421026 45978
rect 421094 45922 421150 45978
rect 421218 45922 421274 45978
rect 421342 45922 421398 45978
rect 420970 28294 421026 28350
rect 421094 28294 421150 28350
rect 421218 28294 421274 28350
rect 421342 28294 421398 28350
rect 420970 28170 421026 28226
rect 421094 28170 421150 28226
rect 421218 28170 421274 28226
rect 421342 28170 421398 28226
rect 420970 28046 421026 28102
rect 421094 28046 421150 28102
rect 421218 28046 421274 28102
rect 421342 28046 421398 28102
rect 420970 27922 421026 27978
rect 421094 27922 421150 27978
rect 421218 27922 421274 27978
rect 421342 27922 421398 27978
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 58294 435306 58350
rect 435374 58294 435430 58350
rect 435498 58294 435554 58350
rect 435622 58294 435678 58350
rect 435250 58170 435306 58226
rect 435374 58170 435430 58226
rect 435498 58170 435554 58226
rect 435622 58170 435678 58226
rect 435250 58046 435306 58102
rect 435374 58046 435430 58102
rect 435498 58046 435554 58102
rect 435622 58046 435678 58102
rect 435250 57922 435306 57978
rect 435374 57922 435430 57978
rect 435498 57922 435554 57978
rect 435622 57922 435678 57978
rect 435250 40294 435306 40350
rect 435374 40294 435430 40350
rect 435498 40294 435554 40350
rect 435622 40294 435678 40350
rect 435250 40170 435306 40226
rect 435374 40170 435430 40226
rect 435498 40170 435554 40226
rect 435622 40170 435678 40226
rect 435250 40046 435306 40102
rect 435374 40046 435430 40102
rect 435498 40046 435554 40102
rect 435622 40046 435678 40102
rect 435250 39922 435306 39978
rect 435374 39922 435430 39978
rect 435498 39922 435554 39978
rect 435622 39922 435678 39978
rect 435250 22294 435306 22350
rect 435374 22294 435430 22350
rect 435498 22294 435554 22350
rect 435622 22294 435678 22350
rect 435250 22170 435306 22226
rect 435374 22170 435430 22226
rect 435498 22170 435554 22226
rect 435622 22170 435678 22226
rect 435250 22046 435306 22102
rect 435374 22046 435430 22102
rect 435498 22046 435554 22102
rect 435622 22046 435678 22102
rect 435250 21922 435306 21978
rect 435374 21922 435430 21978
rect 435498 21922 435554 21978
rect 435622 21922 435678 21978
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 438970 514294 439026 514350
rect 439094 514294 439150 514350
rect 439218 514294 439274 514350
rect 439342 514294 439398 514350
rect 438970 514170 439026 514226
rect 439094 514170 439150 514226
rect 439218 514170 439274 514226
rect 439342 514170 439398 514226
rect 438970 514046 439026 514102
rect 439094 514046 439150 514102
rect 439218 514046 439274 514102
rect 439342 514046 439398 514102
rect 438970 513922 439026 513978
rect 439094 513922 439150 513978
rect 439218 513922 439274 513978
rect 439342 513922 439398 513978
rect 438970 496294 439026 496350
rect 439094 496294 439150 496350
rect 439218 496294 439274 496350
rect 439342 496294 439398 496350
rect 438970 496170 439026 496226
rect 439094 496170 439150 496226
rect 439218 496170 439274 496226
rect 439342 496170 439398 496226
rect 438970 496046 439026 496102
rect 439094 496046 439150 496102
rect 439218 496046 439274 496102
rect 439342 496046 439398 496102
rect 438970 495922 439026 495978
rect 439094 495922 439150 495978
rect 439218 495922 439274 495978
rect 439342 495922 439398 495978
rect 438970 478294 439026 478350
rect 439094 478294 439150 478350
rect 439218 478294 439274 478350
rect 439342 478294 439398 478350
rect 438970 478170 439026 478226
rect 439094 478170 439150 478226
rect 439218 478170 439274 478226
rect 439342 478170 439398 478226
rect 438970 478046 439026 478102
rect 439094 478046 439150 478102
rect 439218 478046 439274 478102
rect 439342 478046 439398 478102
rect 438970 477922 439026 477978
rect 439094 477922 439150 477978
rect 439218 477922 439274 477978
rect 439342 477922 439398 477978
rect 438970 460294 439026 460350
rect 439094 460294 439150 460350
rect 439218 460294 439274 460350
rect 439342 460294 439398 460350
rect 438970 460170 439026 460226
rect 439094 460170 439150 460226
rect 439218 460170 439274 460226
rect 439342 460170 439398 460226
rect 438970 460046 439026 460102
rect 439094 460046 439150 460102
rect 439218 460046 439274 460102
rect 439342 460046 439398 460102
rect 438970 459922 439026 459978
rect 439094 459922 439150 459978
rect 439218 459922 439274 459978
rect 439342 459922 439398 459978
rect 438970 442294 439026 442350
rect 439094 442294 439150 442350
rect 439218 442294 439274 442350
rect 439342 442294 439398 442350
rect 438970 442170 439026 442226
rect 439094 442170 439150 442226
rect 439218 442170 439274 442226
rect 439342 442170 439398 442226
rect 438970 442046 439026 442102
rect 439094 442046 439150 442102
rect 439218 442046 439274 442102
rect 439342 442046 439398 442102
rect 438970 441922 439026 441978
rect 439094 441922 439150 441978
rect 439218 441922 439274 441978
rect 439342 441922 439398 441978
rect 438970 424294 439026 424350
rect 439094 424294 439150 424350
rect 439218 424294 439274 424350
rect 439342 424294 439398 424350
rect 438970 424170 439026 424226
rect 439094 424170 439150 424226
rect 439218 424170 439274 424226
rect 439342 424170 439398 424226
rect 438970 424046 439026 424102
rect 439094 424046 439150 424102
rect 439218 424046 439274 424102
rect 439342 424046 439398 424102
rect 438970 423922 439026 423978
rect 439094 423922 439150 423978
rect 439218 423922 439274 423978
rect 439342 423922 439398 423978
rect 438970 406294 439026 406350
rect 439094 406294 439150 406350
rect 439218 406294 439274 406350
rect 439342 406294 439398 406350
rect 438970 406170 439026 406226
rect 439094 406170 439150 406226
rect 439218 406170 439274 406226
rect 439342 406170 439398 406226
rect 438970 406046 439026 406102
rect 439094 406046 439150 406102
rect 439218 406046 439274 406102
rect 439342 406046 439398 406102
rect 438970 405922 439026 405978
rect 439094 405922 439150 405978
rect 439218 405922 439274 405978
rect 439342 405922 439398 405978
rect 438970 388294 439026 388350
rect 439094 388294 439150 388350
rect 439218 388294 439274 388350
rect 439342 388294 439398 388350
rect 438970 388170 439026 388226
rect 439094 388170 439150 388226
rect 439218 388170 439274 388226
rect 439342 388170 439398 388226
rect 438970 388046 439026 388102
rect 439094 388046 439150 388102
rect 439218 388046 439274 388102
rect 439342 388046 439398 388102
rect 438970 387922 439026 387978
rect 439094 387922 439150 387978
rect 439218 387922 439274 387978
rect 439342 387922 439398 387978
rect 438970 370294 439026 370350
rect 439094 370294 439150 370350
rect 439218 370294 439274 370350
rect 439342 370294 439398 370350
rect 438970 370170 439026 370226
rect 439094 370170 439150 370226
rect 439218 370170 439274 370226
rect 439342 370170 439398 370226
rect 438970 370046 439026 370102
rect 439094 370046 439150 370102
rect 439218 370046 439274 370102
rect 439342 370046 439398 370102
rect 438970 369922 439026 369978
rect 439094 369922 439150 369978
rect 439218 369922 439274 369978
rect 439342 369922 439398 369978
rect 438970 352294 439026 352350
rect 439094 352294 439150 352350
rect 439218 352294 439274 352350
rect 439342 352294 439398 352350
rect 438970 352170 439026 352226
rect 439094 352170 439150 352226
rect 439218 352170 439274 352226
rect 439342 352170 439398 352226
rect 438970 352046 439026 352102
rect 439094 352046 439150 352102
rect 439218 352046 439274 352102
rect 439342 352046 439398 352102
rect 438970 351922 439026 351978
rect 439094 351922 439150 351978
rect 439218 351922 439274 351978
rect 439342 351922 439398 351978
rect 438970 334294 439026 334350
rect 439094 334294 439150 334350
rect 439218 334294 439274 334350
rect 439342 334294 439398 334350
rect 438970 334170 439026 334226
rect 439094 334170 439150 334226
rect 439218 334170 439274 334226
rect 439342 334170 439398 334226
rect 438970 334046 439026 334102
rect 439094 334046 439150 334102
rect 439218 334046 439274 334102
rect 439342 334046 439398 334102
rect 438970 333922 439026 333978
rect 439094 333922 439150 333978
rect 439218 333922 439274 333978
rect 439342 333922 439398 333978
rect 438970 316294 439026 316350
rect 439094 316294 439150 316350
rect 439218 316294 439274 316350
rect 439342 316294 439398 316350
rect 438970 316170 439026 316226
rect 439094 316170 439150 316226
rect 439218 316170 439274 316226
rect 439342 316170 439398 316226
rect 438970 316046 439026 316102
rect 439094 316046 439150 316102
rect 439218 316046 439274 316102
rect 439342 316046 439398 316102
rect 438970 315922 439026 315978
rect 439094 315922 439150 315978
rect 439218 315922 439274 315978
rect 439342 315922 439398 315978
rect 438970 298294 439026 298350
rect 439094 298294 439150 298350
rect 439218 298294 439274 298350
rect 439342 298294 439398 298350
rect 438970 298170 439026 298226
rect 439094 298170 439150 298226
rect 439218 298170 439274 298226
rect 439342 298170 439398 298226
rect 438970 298046 439026 298102
rect 439094 298046 439150 298102
rect 439218 298046 439274 298102
rect 439342 298046 439398 298102
rect 438970 297922 439026 297978
rect 439094 297922 439150 297978
rect 439218 297922 439274 297978
rect 439342 297922 439398 297978
rect 438970 280294 439026 280350
rect 439094 280294 439150 280350
rect 439218 280294 439274 280350
rect 439342 280294 439398 280350
rect 438970 280170 439026 280226
rect 439094 280170 439150 280226
rect 439218 280170 439274 280226
rect 439342 280170 439398 280226
rect 438970 280046 439026 280102
rect 439094 280046 439150 280102
rect 439218 280046 439274 280102
rect 439342 280046 439398 280102
rect 438970 279922 439026 279978
rect 439094 279922 439150 279978
rect 439218 279922 439274 279978
rect 439342 279922 439398 279978
rect 438970 262294 439026 262350
rect 439094 262294 439150 262350
rect 439218 262294 439274 262350
rect 439342 262294 439398 262350
rect 438970 262170 439026 262226
rect 439094 262170 439150 262226
rect 439218 262170 439274 262226
rect 439342 262170 439398 262226
rect 438970 262046 439026 262102
rect 439094 262046 439150 262102
rect 439218 262046 439274 262102
rect 439342 262046 439398 262102
rect 438970 261922 439026 261978
rect 439094 261922 439150 261978
rect 439218 261922 439274 261978
rect 439342 261922 439398 261978
rect 438970 244294 439026 244350
rect 439094 244294 439150 244350
rect 439218 244294 439274 244350
rect 439342 244294 439398 244350
rect 438970 244170 439026 244226
rect 439094 244170 439150 244226
rect 439218 244170 439274 244226
rect 439342 244170 439398 244226
rect 438970 244046 439026 244102
rect 439094 244046 439150 244102
rect 439218 244046 439274 244102
rect 439342 244046 439398 244102
rect 438970 243922 439026 243978
rect 439094 243922 439150 243978
rect 439218 243922 439274 243978
rect 439342 243922 439398 243978
rect 438970 226294 439026 226350
rect 439094 226294 439150 226350
rect 439218 226294 439274 226350
rect 439342 226294 439398 226350
rect 438970 226170 439026 226226
rect 439094 226170 439150 226226
rect 439218 226170 439274 226226
rect 439342 226170 439398 226226
rect 438970 226046 439026 226102
rect 439094 226046 439150 226102
rect 439218 226046 439274 226102
rect 439342 226046 439398 226102
rect 438970 225922 439026 225978
rect 439094 225922 439150 225978
rect 439218 225922 439274 225978
rect 439342 225922 439398 225978
rect 438970 208294 439026 208350
rect 439094 208294 439150 208350
rect 439218 208294 439274 208350
rect 439342 208294 439398 208350
rect 438970 208170 439026 208226
rect 439094 208170 439150 208226
rect 439218 208170 439274 208226
rect 439342 208170 439398 208226
rect 438970 208046 439026 208102
rect 439094 208046 439150 208102
rect 439218 208046 439274 208102
rect 439342 208046 439398 208102
rect 438970 207922 439026 207978
rect 439094 207922 439150 207978
rect 439218 207922 439274 207978
rect 439342 207922 439398 207978
rect 438970 190294 439026 190350
rect 439094 190294 439150 190350
rect 439218 190294 439274 190350
rect 439342 190294 439398 190350
rect 438970 190170 439026 190226
rect 439094 190170 439150 190226
rect 439218 190170 439274 190226
rect 439342 190170 439398 190226
rect 438970 190046 439026 190102
rect 439094 190046 439150 190102
rect 439218 190046 439274 190102
rect 439342 190046 439398 190102
rect 438970 189922 439026 189978
rect 439094 189922 439150 189978
rect 439218 189922 439274 189978
rect 439342 189922 439398 189978
rect 438970 172294 439026 172350
rect 439094 172294 439150 172350
rect 439218 172294 439274 172350
rect 439342 172294 439398 172350
rect 438970 172170 439026 172226
rect 439094 172170 439150 172226
rect 439218 172170 439274 172226
rect 439342 172170 439398 172226
rect 438970 172046 439026 172102
rect 439094 172046 439150 172102
rect 439218 172046 439274 172102
rect 439342 172046 439398 172102
rect 438970 171922 439026 171978
rect 439094 171922 439150 171978
rect 439218 171922 439274 171978
rect 439342 171922 439398 171978
rect 438970 154294 439026 154350
rect 439094 154294 439150 154350
rect 439218 154294 439274 154350
rect 439342 154294 439398 154350
rect 438970 154170 439026 154226
rect 439094 154170 439150 154226
rect 439218 154170 439274 154226
rect 439342 154170 439398 154226
rect 438970 154046 439026 154102
rect 439094 154046 439150 154102
rect 439218 154046 439274 154102
rect 439342 154046 439398 154102
rect 438970 153922 439026 153978
rect 439094 153922 439150 153978
rect 439218 153922 439274 153978
rect 439342 153922 439398 153978
rect 438970 136294 439026 136350
rect 439094 136294 439150 136350
rect 439218 136294 439274 136350
rect 439342 136294 439398 136350
rect 438970 136170 439026 136226
rect 439094 136170 439150 136226
rect 439218 136170 439274 136226
rect 439342 136170 439398 136226
rect 438970 136046 439026 136102
rect 439094 136046 439150 136102
rect 439218 136046 439274 136102
rect 439342 136046 439398 136102
rect 438970 135922 439026 135978
rect 439094 135922 439150 135978
rect 439218 135922 439274 135978
rect 439342 135922 439398 135978
rect 438970 118294 439026 118350
rect 439094 118294 439150 118350
rect 439218 118294 439274 118350
rect 439342 118294 439398 118350
rect 438970 118170 439026 118226
rect 439094 118170 439150 118226
rect 439218 118170 439274 118226
rect 439342 118170 439398 118226
rect 438970 118046 439026 118102
rect 439094 118046 439150 118102
rect 439218 118046 439274 118102
rect 439342 118046 439398 118102
rect 438970 117922 439026 117978
rect 439094 117922 439150 117978
rect 439218 117922 439274 117978
rect 439342 117922 439398 117978
rect 438970 100294 439026 100350
rect 439094 100294 439150 100350
rect 439218 100294 439274 100350
rect 439342 100294 439398 100350
rect 438970 100170 439026 100226
rect 439094 100170 439150 100226
rect 439218 100170 439274 100226
rect 439342 100170 439398 100226
rect 438970 100046 439026 100102
rect 439094 100046 439150 100102
rect 439218 100046 439274 100102
rect 439342 100046 439398 100102
rect 438970 99922 439026 99978
rect 439094 99922 439150 99978
rect 439218 99922 439274 99978
rect 439342 99922 439398 99978
rect 438970 82294 439026 82350
rect 439094 82294 439150 82350
rect 439218 82294 439274 82350
rect 439342 82294 439398 82350
rect 438970 82170 439026 82226
rect 439094 82170 439150 82226
rect 439218 82170 439274 82226
rect 439342 82170 439398 82226
rect 438970 82046 439026 82102
rect 439094 82046 439150 82102
rect 439218 82046 439274 82102
rect 439342 82046 439398 82102
rect 438970 81922 439026 81978
rect 439094 81922 439150 81978
rect 439218 81922 439274 81978
rect 439342 81922 439398 81978
rect 438970 64294 439026 64350
rect 439094 64294 439150 64350
rect 439218 64294 439274 64350
rect 439342 64294 439398 64350
rect 438970 64170 439026 64226
rect 439094 64170 439150 64226
rect 439218 64170 439274 64226
rect 439342 64170 439398 64226
rect 438970 64046 439026 64102
rect 439094 64046 439150 64102
rect 439218 64046 439274 64102
rect 439342 64046 439398 64102
rect 438970 63922 439026 63978
rect 439094 63922 439150 63978
rect 439218 63922 439274 63978
rect 439342 63922 439398 63978
rect 438970 46294 439026 46350
rect 439094 46294 439150 46350
rect 439218 46294 439274 46350
rect 439342 46294 439398 46350
rect 438970 46170 439026 46226
rect 439094 46170 439150 46226
rect 439218 46170 439274 46226
rect 439342 46170 439398 46226
rect 438970 46046 439026 46102
rect 439094 46046 439150 46102
rect 439218 46046 439274 46102
rect 439342 46046 439398 46102
rect 438970 45922 439026 45978
rect 439094 45922 439150 45978
rect 439218 45922 439274 45978
rect 439342 45922 439398 45978
rect 438970 28294 439026 28350
rect 439094 28294 439150 28350
rect 439218 28294 439274 28350
rect 439342 28294 439398 28350
rect 438970 28170 439026 28226
rect 439094 28170 439150 28226
rect 439218 28170 439274 28226
rect 439342 28170 439398 28226
rect 438970 28046 439026 28102
rect 439094 28046 439150 28102
rect 439218 28046 439274 28102
rect 439342 28046 439398 28102
rect 438970 27922 439026 27978
rect 439094 27922 439150 27978
rect 439218 27922 439274 27978
rect 439342 27922 439398 27978
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 453250 526294 453306 526350
rect 453374 526294 453430 526350
rect 453498 526294 453554 526350
rect 453622 526294 453678 526350
rect 453250 526170 453306 526226
rect 453374 526170 453430 526226
rect 453498 526170 453554 526226
rect 453622 526170 453678 526226
rect 453250 526046 453306 526102
rect 453374 526046 453430 526102
rect 453498 526046 453554 526102
rect 453622 526046 453678 526102
rect 453250 525922 453306 525978
rect 453374 525922 453430 525978
rect 453498 525922 453554 525978
rect 453622 525922 453678 525978
rect 453250 508294 453306 508350
rect 453374 508294 453430 508350
rect 453498 508294 453554 508350
rect 453622 508294 453678 508350
rect 453250 508170 453306 508226
rect 453374 508170 453430 508226
rect 453498 508170 453554 508226
rect 453622 508170 453678 508226
rect 453250 508046 453306 508102
rect 453374 508046 453430 508102
rect 453498 508046 453554 508102
rect 453622 508046 453678 508102
rect 453250 507922 453306 507978
rect 453374 507922 453430 507978
rect 453498 507922 453554 507978
rect 453622 507922 453678 507978
rect 453250 490294 453306 490350
rect 453374 490294 453430 490350
rect 453498 490294 453554 490350
rect 453622 490294 453678 490350
rect 453250 490170 453306 490226
rect 453374 490170 453430 490226
rect 453498 490170 453554 490226
rect 453622 490170 453678 490226
rect 453250 490046 453306 490102
rect 453374 490046 453430 490102
rect 453498 490046 453554 490102
rect 453622 490046 453678 490102
rect 453250 489922 453306 489978
rect 453374 489922 453430 489978
rect 453498 489922 453554 489978
rect 453622 489922 453678 489978
rect 453250 472294 453306 472350
rect 453374 472294 453430 472350
rect 453498 472294 453554 472350
rect 453622 472294 453678 472350
rect 453250 472170 453306 472226
rect 453374 472170 453430 472226
rect 453498 472170 453554 472226
rect 453622 472170 453678 472226
rect 453250 472046 453306 472102
rect 453374 472046 453430 472102
rect 453498 472046 453554 472102
rect 453622 472046 453678 472102
rect 453250 471922 453306 471978
rect 453374 471922 453430 471978
rect 453498 471922 453554 471978
rect 453622 471922 453678 471978
rect 453250 454294 453306 454350
rect 453374 454294 453430 454350
rect 453498 454294 453554 454350
rect 453622 454294 453678 454350
rect 453250 454170 453306 454226
rect 453374 454170 453430 454226
rect 453498 454170 453554 454226
rect 453622 454170 453678 454226
rect 453250 454046 453306 454102
rect 453374 454046 453430 454102
rect 453498 454046 453554 454102
rect 453622 454046 453678 454102
rect 453250 453922 453306 453978
rect 453374 453922 453430 453978
rect 453498 453922 453554 453978
rect 453622 453922 453678 453978
rect 453250 436294 453306 436350
rect 453374 436294 453430 436350
rect 453498 436294 453554 436350
rect 453622 436294 453678 436350
rect 453250 436170 453306 436226
rect 453374 436170 453430 436226
rect 453498 436170 453554 436226
rect 453622 436170 453678 436226
rect 453250 436046 453306 436102
rect 453374 436046 453430 436102
rect 453498 436046 453554 436102
rect 453622 436046 453678 436102
rect 453250 435922 453306 435978
rect 453374 435922 453430 435978
rect 453498 435922 453554 435978
rect 453622 435922 453678 435978
rect 453250 418294 453306 418350
rect 453374 418294 453430 418350
rect 453498 418294 453554 418350
rect 453622 418294 453678 418350
rect 453250 418170 453306 418226
rect 453374 418170 453430 418226
rect 453498 418170 453554 418226
rect 453622 418170 453678 418226
rect 453250 418046 453306 418102
rect 453374 418046 453430 418102
rect 453498 418046 453554 418102
rect 453622 418046 453678 418102
rect 453250 417922 453306 417978
rect 453374 417922 453430 417978
rect 453498 417922 453554 417978
rect 453622 417922 453678 417978
rect 453250 400294 453306 400350
rect 453374 400294 453430 400350
rect 453498 400294 453554 400350
rect 453622 400294 453678 400350
rect 453250 400170 453306 400226
rect 453374 400170 453430 400226
rect 453498 400170 453554 400226
rect 453622 400170 453678 400226
rect 453250 400046 453306 400102
rect 453374 400046 453430 400102
rect 453498 400046 453554 400102
rect 453622 400046 453678 400102
rect 453250 399922 453306 399978
rect 453374 399922 453430 399978
rect 453498 399922 453554 399978
rect 453622 399922 453678 399978
rect 453250 382294 453306 382350
rect 453374 382294 453430 382350
rect 453498 382294 453554 382350
rect 453622 382294 453678 382350
rect 453250 382170 453306 382226
rect 453374 382170 453430 382226
rect 453498 382170 453554 382226
rect 453622 382170 453678 382226
rect 453250 382046 453306 382102
rect 453374 382046 453430 382102
rect 453498 382046 453554 382102
rect 453622 382046 453678 382102
rect 453250 381922 453306 381978
rect 453374 381922 453430 381978
rect 453498 381922 453554 381978
rect 453622 381922 453678 381978
rect 453250 364294 453306 364350
rect 453374 364294 453430 364350
rect 453498 364294 453554 364350
rect 453622 364294 453678 364350
rect 453250 364170 453306 364226
rect 453374 364170 453430 364226
rect 453498 364170 453554 364226
rect 453622 364170 453678 364226
rect 453250 364046 453306 364102
rect 453374 364046 453430 364102
rect 453498 364046 453554 364102
rect 453622 364046 453678 364102
rect 453250 363922 453306 363978
rect 453374 363922 453430 363978
rect 453498 363922 453554 363978
rect 453622 363922 453678 363978
rect 453250 346294 453306 346350
rect 453374 346294 453430 346350
rect 453498 346294 453554 346350
rect 453622 346294 453678 346350
rect 453250 346170 453306 346226
rect 453374 346170 453430 346226
rect 453498 346170 453554 346226
rect 453622 346170 453678 346226
rect 453250 346046 453306 346102
rect 453374 346046 453430 346102
rect 453498 346046 453554 346102
rect 453622 346046 453678 346102
rect 453250 345922 453306 345978
rect 453374 345922 453430 345978
rect 453498 345922 453554 345978
rect 453622 345922 453678 345978
rect 453250 328294 453306 328350
rect 453374 328294 453430 328350
rect 453498 328294 453554 328350
rect 453622 328294 453678 328350
rect 453250 328170 453306 328226
rect 453374 328170 453430 328226
rect 453498 328170 453554 328226
rect 453622 328170 453678 328226
rect 453250 328046 453306 328102
rect 453374 328046 453430 328102
rect 453498 328046 453554 328102
rect 453622 328046 453678 328102
rect 453250 327922 453306 327978
rect 453374 327922 453430 327978
rect 453498 327922 453554 327978
rect 453622 327922 453678 327978
rect 453250 310294 453306 310350
rect 453374 310294 453430 310350
rect 453498 310294 453554 310350
rect 453622 310294 453678 310350
rect 453250 310170 453306 310226
rect 453374 310170 453430 310226
rect 453498 310170 453554 310226
rect 453622 310170 453678 310226
rect 453250 310046 453306 310102
rect 453374 310046 453430 310102
rect 453498 310046 453554 310102
rect 453622 310046 453678 310102
rect 453250 309922 453306 309978
rect 453374 309922 453430 309978
rect 453498 309922 453554 309978
rect 453622 309922 453678 309978
rect 453250 292294 453306 292350
rect 453374 292294 453430 292350
rect 453498 292294 453554 292350
rect 453622 292294 453678 292350
rect 453250 292170 453306 292226
rect 453374 292170 453430 292226
rect 453498 292170 453554 292226
rect 453622 292170 453678 292226
rect 453250 292046 453306 292102
rect 453374 292046 453430 292102
rect 453498 292046 453554 292102
rect 453622 292046 453678 292102
rect 453250 291922 453306 291978
rect 453374 291922 453430 291978
rect 453498 291922 453554 291978
rect 453622 291922 453678 291978
rect 453250 274294 453306 274350
rect 453374 274294 453430 274350
rect 453498 274294 453554 274350
rect 453622 274294 453678 274350
rect 453250 274170 453306 274226
rect 453374 274170 453430 274226
rect 453498 274170 453554 274226
rect 453622 274170 453678 274226
rect 453250 274046 453306 274102
rect 453374 274046 453430 274102
rect 453498 274046 453554 274102
rect 453622 274046 453678 274102
rect 453250 273922 453306 273978
rect 453374 273922 453430 273978
rect 453498 273922 453554 273978
rect 453622 273922 453678 273978
rect 453250 256294 453306 256350
rect 453374 256294 453430 256350
rect 453498 256294 453554 256350
rect 453622 256294 453678 256350
rect 453250 256170 453306 256226
rect 453374 256170 453430 256226
rect 453498 256170 453554 256226
rect 453622 256170 453678 256226
rect 453250 256046 453306 256102
rect 453374 256046 453430 256102
rect 453498 256046 453554 256102
rect 453622 256046 453678 256102
rect 453250 255922 453306 255978
rect 453374 255922 453430 255978
rect 453498 255922 453554 255978
rect 453622 255922 453678 255978
rect 453250 238294 453306 238350
rect 453374 238294 453430 238350
rect 453498 238294 453554 238350
rect 453622 238294 453678 238350
rect 453250 238170 453306 238226
rect 453374 238170 453430 238226
rect 453498 238170 453554 238226
rect 453622 238170 453678 238226
rect 453250 238046 453306 238102
rect 453374 238046 453430 238102
rect 453498 238046 453554 238102
rect 453622 238046 453678 238102
rect 453250 237922 453306 237978
rect 453374 237922 453430 237978
rect 453498 237922 453554 237978
rect 453622 237922 453678 237978
rect 453250 220294 453306 220350
rect 453374 220294 453430 220350
rect 453498 220294 453554 220350
rect 453622 220294 453678 220350
rect 453250 220170 453306 220226
rect 453374 220170 453430 220226
rect 453498 220170 453554 220226
rect 453622 220170 453678 220226
rect 453250 220046 453306 220102
rect 453374 220046 453430 220102
rect 453498 220046 453554 220102
rect 453622 220046 453678 220102
rect 453250 219922 453306 219978
rect 453374 219922 453430 219978
rect 453498 219922 453554 219978
rect 453622 219922 453678 219978
rect 453250 202294 453306 202350
rect 453374 202294 453430 202350
rect 453498 202294 453554 202350
rect 453622 202294 453678 202350
rect 453250 202170 453306 202226
rect 453374 202170 453430 202226
rect 453498 202170 453554 202226
rect 453622 202170 453678 202226
rect 453250 202046 453306 202102
rect 453374 202046 453430 202102
rect 453498 202046 453554 202102
rect 453622 202046 453678 202102
rect 453250 201922 453306 201978
rect 453374 201922 453430 201978
rect 453498 201922 453554 201978
rect 453622 201922 453678 201978
rect 453250 184294 453306 184350
rect 453374 184294 453430 184350
rect 453498 184294 453554 184350
rect 453622 184294 453678 184350
rect 453250 184170 453306 184226
rect 453374 184170 453430 184226
rect 453498 184170 453554 184226
rect 453622 184170 453678 184226
rect 453250 184046 453306 184102
rect 453374 184046 453430 184102
rect 453498 184046 453554 184102
rect 453622 184046 453678 184102
rect 453250 183922 453306 183978
rect 453374 183922 453430 183978
rect 453498 183922 453554 183978
rect 453622 183922 453678 183978
rect 453250 166294 453306 166350
rect 453374 166294 453430 166350
rect 453498 166294 453554 166350
rect 453622 166294 453678 166350
rect 453250 166170 453306 166226
rect 453374 166170 453430 166226
rect 453498 166170 453554 166226
rect 453622 166170 453678 166226
rect 453250 166046 453306 166102
rect 453374 166046 453430 166102
rect 453498 166046 453554 166102
rect 453622 166046 453678 166102
rect 453250 165922 453306 165978
rect 453374 165922 453430 165978
rect 453498 165922 453554 165978
rect 453622 165922 453678 165978
rect 453250 148294 453306 148350
rect 453374 148294 453430 148350
rect 453498 148294 453554 148350
rect 453622 148294 453678 148350
rect 453250 148170 453306 148226
rect 453374 148170 453430 148226
rect 453498 148170 453554 148226
rect 453622 148170 453678 148226
rect 453250 148046 453306 148102
rect 453374 148046 453430 148102
rect 453498 148046 453554 148102
rect 453622 148046 453678 148102
rect 453250 147922 453306 147978
rect 453374 147922 453430 147978
rect 453498 147922 453554 147978
rect 453622 147922 453678 147978
rect 453250 130294 453306 130350
rect 453374 130294 453430 130350
rect 453498 130294 453554 130350
rect 453622 130294 453678 130350
rect 453250 130170 453306 130226
rect 453374 130170 453430 130226
rect 453498 130170 453554 130226
rect 453622 130170 453678 130226
rect 453250 130046 453306 130102
rect 453374 130046 453430 130102
rect 453498 130046 453554 130102
rect 453622 130046 453678 130102
rect 453250 129922 453306 129978
rect 453374 129922 453430 129978
rect 453498 129922 453554 129978
rect 453622 129922 453678 129978
rect 453250 112294 453306 112350
rect 453374 112294 453430 112350
rect 453498 112294 453554 112350
rect 453622 112294 453678 112350
rect 453250 112170 453306 112226
rect 453374 112170 453430 112226
rect 453498 112170 453554 112226
rect 453622 112170 453678 112226
rect 453250 112046 453306 112102
rect 453374 112046 453430 112102
rect 453498 112046 453554 112102
rect 453622 112046 453678 112102
rect 453250 111922 453306 111978
rect 453374 111922 453430 111978
rect 453498 111922 453554 111978
rect 453622 111922 453678 111978
rect 453250 94294 453306 94350
rect 453374 94294 453430 94350
rect 453498 94294 453554 94350
rect 453622 94294 453678 94350
rect 453250 94170 453306 94226
rect 453374 94170 453430 94226
rect 453498 94170 453554 94226
rect 453622 94170 453678 94226
rect 453250 94046 453306 94102
rect 453374 94046 453430 94102
rect 453498 94046 453554 94102
rect 453622 94046 453678 94102
rect 453250 93922 453306 93978
rect 453374 93922 453430 93978
rect 453498 93922 453554 93978
rect 453622 93922 453678 93978
rect 453250 76294 453306 76350
rect 453374 76294 453430 76350
rect 453498 76294 453554 76350
rect 453622 76294 453678 76350
rect 453250 76170 453306 76226
rect 453374 76170 453430 76226
rect 453498 76170 453554 76226
rect 453622 76170 453678 76226
rect 453250 76046 453306 76102
rect 453374 76046 453430 76102
rect 453498 76046 453554 76102
rect 453622 76046 453678 76102
rect 453250 75922 453306 75978
rect 453374 75922 453430 75978
rect 453498 75922 453554 75978
rect 453622 75922 453678 75978
rect 453250 58294 453306 58350
rect 453374 58294 453430 58350
rect 453498 58294 453554 58350
rect 453622 58294 453678 58350
rect 453250 58170 453306 58226
rect 453374 58170 453430 58226
rect 453498 58170 453554 58226
rect 453622 58170 453678 58226
rect 453250 58046 453306 58102
rect 453374 58046 453430 58102
rect 453498 58046 453554 58102
rect 453622 58046 453678 58102
rect 453250 57922 453306 57978
rect 453374 57922 453430 57978
rect 453498 57922 453554 57978
rect 453622 57922 453678 57978
rect 453250 40294 453306 40350
rect 453374 40294 453430 40350
rect 453498 40294 453554 40350
rect 453622 40294 453678 40350
rect 453250 40170 453306 40226
rect 453374 40170 453430 40226
rect 453498 40170 453554 40226
rect 453622 40170 453678 40226
rect 453250 40046 453306 40102
rect 453374 40046 453430 40102
rect 453498 40046 453554 40102
rect 453622 40046 453678 40102
rect 453250 39922 453306 39978
rect 453374 39922 453430 39978
rect 453498 39922 453554 39978
rect 453622 39922 453678 39978
rect 453250 22294 453306 22350
rect 453374 22294 453430 22350
rect 453498 22294 453554 22350
rect 453622 22294 453678 22350
rect 453250 22170 453306 22226
rect 453374 22170 453430 22226
rect 453498 22170 453554 22226
rect 453622 22170 453678 22226
rect 453250 22046 453306 22102
rect 453374 22046 453430 22102
rect 453498 22046 453554 22102
rect 453622 22046 453678 22102
rect 453250 21922 453306 21978
rect 453374 21922 453430 21978
rect 453498 21922 453554 21978
rect 453622 21922 453678 21978
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 456970 514294 457026 514350
rect 457094 514294 457150 514350
rect 457218 514294 457274 514350
rect 457342 514294 457398 514350
rect 456970 514170 457026 514226
rect 457094 514170 457150 514226
rect 457218 514170 457274 514226
rect 457342 514170 457398 514226
rect 456970 514046 457026 514102
rect 457094 514046 457150 514102
rect 457218 514046 457274 514102
rect 457342 514046 457398 514102
rect 456970 513922 457026 513978
rect 457094 513922 457150 513978
rect 457218 513922 457274 513978
rect 457342 513922 457398 513978
rect 456970 496294 457026 496350
rect 457094 496294 457150 496350
rect 457218 496294 457274 496350
rect 457342 496294 457398 496350
rect 456970 496170 457026 496226
rect 457094 496170 457150 496226
rect 457218 496170 457274 496226
rect 457342 496170 457398 496226
rect 456970 496046 457026 496102
rect 457094 496046 457150 496102
rect 457218 496046 457274 496102
rect 457342 496046 457398 496102
rect 456970 495922 457026 495978
rect 457094 495922 457150 495978
rect 457218 495922 457274 495978
rect 457342 495922 457398 495978
rect 456970 478294 457026 478350
rect 457094 478294 457150 478350
rect 457218 478294 457274 478350
rect 457342 478294 457398 478350
rect 456970 478170 457026 478226
rect 457094 478170 457150 478226
rect 457218 478170 457274 478226
rect 457342 478170 457398 478226
rect 456970 478046 457026 478102
rect 457094 478046 457150 478102
rect 457218 478046 457274 478102
rect 457342 478046 457398 478102
rect 456970 477922 457026 477978
rect 457094 477922 457150 477978
rect 457218 477922 457274 477978
rect 457342 477922 457398 477978
rect 456970 460294 457026 460350
rect 457094 460294 457150 460350
rect 457218 460294 457274 460350
rect 457342 460294 457398 460350
rect 456970 460170 457026 460226
rect 457094 460170 457150 460226
rect 457218 460170 457274 460226
rect 457342 460170 457398 460226
rect 456970 460046 457026 460102
rect 457094 460046 457150 460102
rect 457218 460046 457274 460102
rect 457342 460046 457398 460102
rect 456970 459922 457026 459978
rect 457094 459922 457150 459978
rect 457218 459922 457274 459978
rect 457342 459922 457398 459978
rect 456970 442294 457026 442350
rect 457094 442294 457150 442350
rect 457218 442294 457274 442350
rect 457342 442294 457398 442350
rect 456970 442170 457026 442226
rect 457094 442170 457150 442226
rect 457218 442170 457274 442226
rect 457342 442170 457398 442226
rect 456970 442046 457026 442102
rect 457094 442046 457150 442102
rect 457218 442046 457274 442102
rect 457342 442046 457398 442102
rect 456970 441922 457026 441978
rect 457094 441922 457150 441978
rect 457218 441922 457274 441978
rect 457342 441922 457398 441978
rect 456970 424294 457026 424350
rect 457094 424294 457150 424350
rect 457218 424294 457274 424350
rect 457342 424294 457398 424350
rect 456970 424170 457026 424226
rect 457094 424170 457150 424226
rect 457218 424170 457274 424226
rect 457342 424170 457398 424226
rect 456970 424046 457026 424102
rect 457094 424046 457150 424102
rect 457218 424046 457274 424102
rect 457342 424046 457398 424102
rect 456970 423922 457026 423978
rect 457094 423922 457150 423978
rect 457218 423922 457274 423978
rect 457342 423922 457398 423978
rect 456970 406294 457026 406350
rect 457094 406294 457150 406350
rect 457218 406294 457274 406350
rect 457342 406294 457398 406350
rect 456970 406170 457026 406226
rect 457094 406170 457150 406226
rect 457218 406170 457274 406226
rect 457342 406170 457398 406226
rect 456970 406046 457026 406102
rect 457094 406046 457150 406102
rect 457218 406046 457274 406102
rect 457342 406046 457398 406102
rect 456970 405922 457026 405978
rect 457094 405922 457150 405978
rect 457218 405922 457274 405978
rect 457342 405922 457398 405978
rect 456970 388294 457026 388350
rect 457094 388294 457150 388350
rect 457218 388294 457274 388350
rect 457342 388294 457398 388350
rect 456970 388170 457026 388226
rect 457094 388170 457150 388226
rect 457218 388170 457274 388226
rect 457342 388170 457398 388226
rect 456970 388046 457026 388102
rect 457094 388046 457150 388102
rect 457218 388046 457274 388102
rect 457342 388046 457398 388102
rect 456970 387922 457026 387978
rect 457094 387922 457150 387978
rect 457218 387922 457274 387978
rect 457342 387922 457398 387978
rect 456970 370294 457026 370350
rect 457094 370294 457150 370350
rect 457218 370294 457274 370350
rect 457342 370294 457398 370350
rect 456970 370170 457026 370226
rect 457094 370170 457150 370226
rect 457218 370170 457274 370226
rect 457342 370170 457398 370226
rect 456970 370046 457026 370102
rect 457094 370046 457150 370102
rect 457218 370046 457274 370102
rect 457342 370046 457398 370102
rect 456970 369922 457026 369978
rect 457094 369922 457150 369978
rect 457218 369922 457274 369978
rect 457342 369922 457398 369978
rect 456970 352294 457026 352350
rect 457094 352294 457150 352350
rect 457218 352294 457274 352350
rect 457342 352294 457398 352350
rect 456970 352170 457026 352226
rect 457094 352170 457150 352226
rect 457218 352170 457274 352226
rect 457342 352170 457398 352226
rect 456970 352046 457026 352102
rect 457094 352046 457150 352102
rect 457218 352046 457274 352102
rect 457342 352046 457398 352102
rect 456970 351922 457026 351978
rect 457094 351922 457150 351978
rect 457218 351922 457274 351978
rect 457342 351922 457398 351978
rect 456970 334294 457026 334350
rect 457094 334294 457150 334350
rect 457218 334294 457274 334350
rect 457342 334294 457398 334350
rect 456970 334170 457026 334226
rect 457094 334170 457150 334226
rect 457218 334170 457274 334226
rect 457342 334170 457398 334226
rect 456970 334046 457026 334102
rect 457094 334046 457150 334102
rect 457218 334046 457274 334102
rect 457342 334046 457398 334102
rect 456970 333922 457026 333978
rect 457094 333922 457150 333978
rect 457218 333922 457274 333978
rect 457342 333922 457398 333978
rect 456970 316294 457026 316350
rect 457094 316294 457150 316350
rect 457218 316294 457274 316350
rect 457342 316294 457398 316350
rect 456970 316170 457026 316226
rect 457094 316170 457150 316226
rect 457218 316170 457274 316226
rect 457342 316170 457398 316226
rect 456970 316046 457026 316102
rect 457094 316046 457150 316102
rect 457218 316046 457274 316102
rect 457342 316046 457398 316102
rect 456970 315922 457026 315978
rect 457094 315922 457150 315978
rect 457218 315922 457274 315978
rect 457342 315922 457398 315978
rect 456970 298294 457026 298350
rect 457094 298294 457150 298350
rect 457218 298294 457274 298350
rect 457342 298294 457398 298350
rect 456970 298170 457026 298226
rect 457094 298170 457150 298226
rect 457218 298170 457274 298226
rect 457342 298170 457398 298226
rect 456970 298046 457026 298102
rect 457094 298046 457150 298102
rect 457218 298046 457274 298102
rect 457342 298046 457398 298102
rect 456970 297922 457026 297978
rect 457094 297922 457150 297978
rect 457218 297922 457274 297978
rect 457342 297922 457398 297978
rect 456970 280294 457026 280350
rect 457094 280294 457150 280350
rect 457218 280294 457274 280350
rect 457342 280294 457398 280350
rect 456970 280170 457026 280226
rect 457094 280170 457150 280226
rect 457218 280170 457274 280226
rect 457342 280170 457398 280226
rect 456970 280046 457026 280102
rect 457094 280046 457150 280102
rect 457218 280046 457274 280102
rect 457342 280046 457398 280102
rect 456970 279922 457026 279978
rect 457094 279922 457150 279978
rect 457218 279922 457274 279978
rect 457342 279922 457398 279978
rect 456970 262294 457026 262350
rect 457094 262294 457150 262350
rect 457218 262294 457274 262350
rect 457342 262294 457398 262350
rect 456970 262170 457026 262226
rect 457094 262170 457150 262226
rect 457218 262170 457274 262226
rect 457342 262170 457398 262226
rect 456970 262046 457026 262102
rect 457094 262046 457150 262102
rect 457218 262046 457274 262102
rect 457342 262046 457398 262102
rect 456970 261922 457026 261978
rect 457094 261922 457150 261978
rect 457218 261922 457274 261978
rect 457342 261922 457398 261978
rect 456970 244294 457026 244350
rect 457094 244294 457150 244350
rect 457218 244294 457274 244350
rect 457342 244294 457398 244350
rect 456970 244170 457026 244226
rect 457094 244170 457150 244226
rect 457218 244170 457274 244226
rect 457342 244170 457398 244226
rect 456970 244046 457026 244102
rect 457094 244046 457150 244102
rect 457218 244046 457274 244102
rect 457342 244046 457398 244102
rect 456970 243922 457026 243978
rect 457094 243922 457150 243978
rect 457218 243922 457274 243978
rect 457342 243922 457398 243978
rect 456970 226294 457026 226350
rect 457094 226294 457150 226350
rect 457218 226294 457274 226350
rect 457342 226294 457398 226350
rect 456970 226170 457026 226226
rect 457094 226170 457150 226226
rect 457218 226170 457274 226226
rect 457342 226170 457398 226226
rect 456970 226046 457026 226102
rect 457094 226046 457150 226102
rect 457218 226046 457274 226102
rect 457342 226046 457398 226102
rect 456970 225922 457026 225978
rect 457094 225922 457150 225978
rect 457218 225922 457274 225978
rect 457342 225922 457398 225978
rect 456970 208294 457026 208350
rect 457094 208294 457150 208350
rect 457218 208294 457274 208350
rect 457342 208294 457398 208350
rect 456970 208170 457026 208226
rect 457094 208170 457150 208226
rect 457218 208170 457274 208226
rect 457342 208170 457398 208226
rect 456970 208046 457026 208102
rect 457094 208046 457150 208102
rect 457218 208046 457274 208102
rect 457342 208046 457398 208102
rect 456970 207922 457026 207978
rect 457094 207922 457150 207978
rect 457218 207922 457274 207978
rect 457342 207922 457398 207978
rect 456970 190294 457026 190350
rect 457094 190294 457150 190350
rect 457218 190294 457274 190350
rect 457342 190294 457398 190350
rect 456970 190170 457026 190226
rect 457094 190170 457150 190226
rect 457218 190170 457274 190226
rect 457342 190170 457398 190226
rect 456970 190046 457026 190102
rect 457094 190046 457150 190102
rect 457218 190046 457274 190102
rect 457342 190046 457398 190102
rect 456970 189922 457026 189978
rect 457094 189922 457150 189978
rect 457218 189922 457274 189978
rect 457342 189922 457398 189978
rect 456970 172294 457026 172350
rect 457094 172294 457150 172350
rect 457218 172294 457274 172350
rect 457342 172294 457398 172350
rect 456970 172170 457026 172226
rect 457094 172170 457150 172226
rect 457218 172170 457274 172226
rect 457342 172170 457398 172226
rect 456970 172046 457026 172102
rect 457094 172046 457150 172102
rect 457218 172046 457274 172102
rect 457342 172046 457398 172102
rect 456970 171922 457026 171978
rect 457094 171922 457150 171978
rect 457218 171922 457274 171978
rect 457342 171922 457398 171978
rect 456970 154294 457026 154350
rect 457094 154294 457150 154350
rect 457218 154294 457274 154350
rect 457342 154294 457398 154350
rect 456970 154170 457026 154226
rect 457094 154170 457150 154226
rect 457218 154170 457274 154226
rect 457342 154170 457398 154226
rect 456970 154046 457026 154102
rect 457094 154046 457150 154102
rect 457218 154046 457274 154102
rect 457342 154046 457398 154102
rect 456970 153922 457026 153978
rect 457094 153922 457150 153978
rect 457218 153922 457274 153978
rect 457342 153922 457398 153978
rect 456970 136294 457026 136350
rect 457094 136294 457150 136350
rect 457218 136294 457274 136350
rect 457342 136294 457398 136350
rect 456970 136170 457026 136226
rect 457094 136170 457150 136226
rect 457218 136170 457274 136226
rect 457342 136170 457398 136226
rect 456970 136046 457026 136102
rect 457094 136046 457150 136102
rect 457218 136046 457274 136102
rect 457342 136046 457398 136102
rect 456970 135922 457026 135978
rect 457094 135922 457150 135978
rect 457218 135922 457274 135978
rect 457342 135922 457398 135978
rect 456970 118294 457026 118350
rect 457094 118294 457150 118350
rect 457218 118294 457274 118350
rect 457342 118294 457398 118350
rect 456970 118170 457026 118226
rect 457094 118170 457150 118226
rect 457218 118170 457274 118226
rect 457342 118170 457398 118226
rect 456970 118046 457026 118102
rect 457094 118046 457150 118102
rect 457218 118046 457274 118102
rect 457342 118046 457398 118102
rect 456970 117922 457026 117978
rect 457094 117922 457150 117978
rect 457218 117922 457274 117978
rect 457342 117922 457398 117978
rect 456970 100294 457026 100350
rect 457094 100294 457150 100350
rect 457218 100294 457274 100350
rect 457342 100294 457398 100350
rect 456970 100170 457026 100226
rect 457094 100170 457150 100226
rect 457218 100170 457274 100226
rect 457342 100170 457398 100226
rect 456970 100046 457026 100102
rect 457094 100046 457150 100102
rect 457218 100046 457274 100102
rect 457342 100046 457398 100102
rect 456970 99922 457026 99978
rect 457094 99922 457150 99978
rect 457218 99922 457274 99978
rect 457342 99922 457398 99978
rect 456970 82294 457026 82350
rect 457094 82294 457150 82350
rect 457218 82294 457274 82350
rect 457342 82294 457398 82350
rect 456970 82170 457026 82226
rect 457094 82170 457150 82226
rect 457218 82170 457274 82226
rect 457342 82170 457398 82226
rect 456970 82046 457026 82102
rect 457094 82046 457150 82102
rect 457218 82046 457274 82102
rect 457342 82046 457398 82102
rect 456970 81922 457026 81978
rect 457094 81922 457150 81978
rect 457218 81922 457274 81978
rect 457342 81922 457398 81978
rect 456970 64294 457026 64350
rect 457094 64294 457150 64350
rect 457218 64294 457274 64350
rect 457342 64294 457398 64350
rect 456970 64170 457026 64226
rect 457094 64170 457150 64226
rect 457218 64170 457274 64226
rect 457342 64170 457398 64226
rect 456970 64046 457026 64102
rect 457094 64046 457150 64102
rect 457218 64046 457274 64102
rect 457342 64046 457398 64102
rect 456970 63922 457026 63978
rect 457094 63922 457150 63978
rect 457218 63922 457274 63978
rect 457342 63922 457398 63978
rect 456970 46294 457026 46350
rect 457094 46294 457150 46350
rect 457218 46294 457274 46350
rect 457342 46294 457398 46350
rect 456970 46170 457026 46226
rect 457094 46170 457150 46226
rect 457218 46170 457274 46226
rect 457342 46170 457398 46226
rect 456970 46046 457026 46102
rect 457094 46046 457150 46102
rect 457218 46046 457274 46102
rect 457342 46046 457398 46102
rect 456970 45922 457026 45978
rect 457094 45922 457150 45978
rect 457218 45922 457274 45978
rect 457342 45922 457398 45978
rect 456970 28294 457026 28350
rect 457094 28294 457150 28350
rect 457218 28294 457274 28350
rect 457342 28294 457398 28350
rect 456970 28170 457026 28226
rect 457094 28170 457150 28226
rect 457218 28170 457274 28226
rect 457342 28170 457398 28226
rect 456970 28046 457026 28102
rect 457094 28046 457150 28102
rect 457218 28046 457274 28102
rect 457342 28046 457398 28102
rect 456970 27922 457026 27978
rect 457094 27922 457150 27978
rect 457218 27922 457274 27978
rect 457342 27922 457398 27978
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 471250 526294 471306 526350
rect 471374 526294 471430 526350
rect 471498 526294 471554 526350
rect 471622 526294 471678 526350
rect 471250 526170 471306 526226
rect 471374 526170 471430 526226
rect 471498 526170 471554 526226
rect 471622 526170 471678 526226
rect 471250 526046 471306 526102
rect 471374 526046 471430 526102
rect 471498 526046 471554 526102
rect 471622 526046 471678 526102
rect 471250 525922 471306 525978
rect 471374 525922 471430 525978
rect 471498 525922 471554 525978
rect 471622 525922 471678 525978
rect 471250 508294 471306 508350
rect 471374 508294 471430 508350
rect 471498 508294 471554 508350
rect 471622 508294 471678 508350
rect 471250 508170 471306 508226
rect 471374 508170 471430 508226
rect 471498 508170 471554 508226
rect 471622 508170 471678 508226
rect 471250 508046 471306 508102
rect 471374 508046 471430 508102
rect 471498 508046 471554 508102
rect 471622 508046 471678 508102
rect 471250 507922 471306 507978
rect 471374 507922 471430 507978
rect 471498 507922 471554 507978
rect 471622 507922 471678 507978
rect 471250 490294 471306 490350
rect 471374 490294 471430 490350
rect 471498 490294 471554 490350
rect 471622 490294 471678 490350
rect 471250 490170 471306 490226
rect 471374 490170 471430 490226
rect 471498 490170 471554 490226
rect 471622 490170 471678 490226
rect 471250 490046 471306 490102
rect 471374 490046 471430 490102
rect 471498 490046 471554 490102
rect 471622 490046 471678 490102
rect 471250 489922 471306 489978
rect 471374 489922 471430 489978
rect 471498 489922 471554 489978
rect 471622 489922 471678 489978
rect 471250 472294 471306 472350
rect 471374 472294 471430 472350
rect 471498 472294 471554 472350
rect 471622 472294 471678 472350
rect 471250 472170 471306 472226
rect 471374 472170 471430 472226
rect 471498 472170 471554 472226
rect 471622 472170 471678 472226
rect 471250 472046 471306 472102
rect 471374 472046 471430 472102
rect 471498 472046 471554 472102
rect 471622 472046 471678 472102
rect 471250 471922 471306 471978
rect 471374 471922 471430 471978
rect 471498 471922 471554 471978
rect 471622 471922 471678 471978
rect 471250 454294 471306 454350
rect 471374 454294 471430 454350
rect 471498 454294 471554 454350
rect 471622 454294 471678 454350
rect 471250 454170 471306 454226
rect 471374 454170 471430 454226
rect 471498 454170 471554 454226
rect 471622 454170 471678 454226
rect 471250 454046 471306 454102
rect 471374 454046 471430 454102
rect 471498 454046 471554 454102
rect 471622 454046 471678 454102
rect 471250 453922 471306 453978
rect 471374 453922 471430 453978
rect 471498 453922 471554 453978
rect 471622 453922 471678 453978
rect 471250 436294 471306 436350
rect 471374 436294 471430 436350
rect 471498 436294 471554 436350
rect 471622 436294 471678 436350
rect 471250 436170 471306 436226
rect 471374 436170 471430 436226
rect 471498 436170 471554 436226
rect 471622 436170 471678 436226
rect 471250 436046 471306 436102
rect 471374 436046 471430 436102
rect 471498 436046 471554 436102
rect 471622 436046 471678 436102
rect 471250 435922 471306 435978
rect 471374 435922 471430 435978
rect 471498 435922 471554 435978
rect 471622 435922 471678 435978
rect 471250 418294 471306 418350
rect 471374 418294 471430 418350
rect 471498 418294 471554 418350
rect 471622 418294 471678 418350
rect 471250 418170 471306 418226
rect 471374 418170 471430 418226
rect 471498 418170 471554 418226
rect 471622 418170 471678 418226
rect 471250 418046 471306 418102
rect 471374 418046 471430 418102
rect 471498 418046 471554 418102
rect 471622 418046 471678 418102
rect 471250 417922 471306 417978
rect 471374 417922 471430 417978
rect 471498 417922 471554 417978
rect 471622 417922 471678 417978
rect 471250 400294 471306 400350
rect 471374 400294 471430 400350
rect 471498 400294 471554 400350
rect 471622 400294 471678 400350
rect 471250 400170 471306 400226
rect 471374 400170 471430 400226
rect 471498 400170 471554 400226
rect 471622 400170 471678 400226
rect 471250 400046 471306 400102
rect 471374 400046 471430 400102
rect 471498 400046 471554 400102
rect 471622 400046 471678 400102
rect 471250 399922 471306 399978
rect 471374 399922 471430 399978
rect 471498 399922 471554 399978
rect 471622 399922 471678 399978
rect 471250 382294 471306 382350
rect 471374 382294 471430 382350
rect 471498 382294 471554 382350
rect 471622 382294 471678 382350
rect 471250 382170 471306 382226
rect 471374 382170 471430 382226
rect 471498 382170 471554 382226
rect 471622 382170 471678 382226
rect 471250 382046 471306 382102
rect 471374 382046 471430 382102
rect 471498 382046 471554 382102
rect 471622 382046 471678 382102
rect 471250 381922 471306 381978
rect 471374 381922 471430 381978
rect 471498 381922 471554 381978
rect 471622 381922 471678 381978
rect 471250 364294 471306 364350
rect 471374 364294 471430 364350
rect 471498 364294 471554 364350
rect 471622 364294 471678 364350
rect 471250 364170 471306 364226
rect 471374 364170 471430 364226
rect 471498 364170 471554 364226
rect 471622 364170 471678 364226
rect 471250 364046 471306 364102
rect 471374 364046 471430 364102
rect 471498 364046 471554 364102
rect 471622 364046 471678 364102
rect 471250 363922 471306 363978
rect 471374 363922 471430 363978
rect 471498 363922 471554 363978
rect 471622 363922 471678 363978
rect 471250 346294 471306 346350
rect 471374 346294 471430 346350
rect 471498 346294 471554 346350
rect 471622 346294 471678 346350
rect 471250 346170 471306 346226
rect 471374 346170 471430 346226
rect 471498 346170 471554 346226
rect 471622 346170 471678 346226
rect 471250 346046 471306 346102
rect 471374 346046 471430 346102
rect 471498 346046 471554 346102
rect 471622 346046 471678 346102
rect 471250 345922 471306 345978
rect 471374 345922 471430 345978
rect 471498 345922 471554 345978
rect 471622 345922 471678 345978
rect 471250 328294 471306 328350
rect 471374 328294 471430 328350
rect 471498 328294 471554 328350
rect 471622 328294 471678 328350
rect 471250 328170 471306 328226
rect 471374 328170 471430 328226
rect 471498 328170 471554 328226
rect 471622 328170 471678 328226
rect 471250 328046 471306 328102
rect 471374 328046 471430 328102
rect 471498 328046 471554 328102
rect 471622 328046 471678 328102
rect 471250 327922 471306 327978
rect 471374 327922 471430 327978
rect 471498 327922 471554 327978
rect 471622 327922 471678 327978
rect 471250 310294 471306 310350
rect 471374 310294 471430 310350
rect 471498 310294 471554 310350
rect 471622 310294 471678 310350
rect 471250 310170 471306 310226
rect 471374 310170 471430 310226
rect 471498 310170 471554 310226
rect 471622 310170 471678 310226
rect 471250 310046 471306 310102
rect 471374 310046 471430 310102
rect 471498 310046 471554 310102
rect 471622 310046 471678 310102
rect 471250 309922 471306 309978
rect 471374 309922 471430 309978
rect 471498 309922 471554 309978
rect 471622 309922 471678 309978
rect 471250 292294 471306 292350
rect 471374 292294 471430 292350
rect 471498 292294 471554 292350
rect 471622 292294 471678 292350
rect 471250 292170 471306 292226
rect 471374 292170 471430 292226
rect 471498 292170 471554 292226
rect 471622 292170 471678 292226
rect 471250 292046 471306 292102
rect 471374 292046 471430 292102
rect 471498 292046 471554 292102
rect 471622 292046 471678 292102
rect 471250 291922 471306 291978
rect 471374 291922 471430 291978
rect 471498 291922 471554 291978
rect 471622 291922 471678 291978
rect 471250 274294 471306 274350
rect 471374 274294 471430 274350
rect 471498 274294 471554 274350
rect 471622 274294 471678 274350
rect 471250 274170 471306 274226
rect 471374 274170 471430 274226
rect 471498 274170 471554 274226
rect 471622 274170 471678 274226
rect 471250 274046 471306 274102
rect 471374 274046 471430 274102
rect 471498 274046 471554 274102
rect 471622 274046 471678 274102
rect 471250 273922 471306 273978
rect 471374 273922 471430 273978
rect 471498 273922 471554 273978
rect 471622 273922 471678 273978
rect 471250 256294 471306 256350
rect 471374 256294 471430 256350
rect 471498 256294 471554 256350
rect 471622 256294 471678 256350
rect 471250 256170 471306 256226
rect 471374 256170 471430 256226
rect 471498 256170 471554 256226
rect 471622 256170 471678 256226
rect 471250 256046 471306 256102
rect 471374 256046 471430 256102
rect 471498 256046 471554 256102
rect 471622 256046 471678 256102
rect 471250 255922 471306 255978
rect 471374 255922 471430 255978
rect 471498 255922 471554 255978
rect 471622 255922 471678 255978
rect 471250 238294 471306 238350
rect 471374 238294 471430 238350
rect 471498 238294 471554 238350
rect 471622 238294 471678 238350
rect 471250 238170 471306 238226
rect 471374 238170 471430 238226
rect 471498 238170 471554 238226
rect 471622 238170 471678 238226
rect 471250 238046 471306 238102
rect 471374 238046 471430 238102
rect 471498 238046 471554 238102
rect 471622 238046 471678 238102
rect 471250 237922 471306 237978
rect 471374 237922 471430 237978
rect 471498 237922 471554 237978
rect 471622 237922 471678 237978
rect 471250 220294 471306 220350
rect 471374 220294 471430 220350
rect 471498 220294 471554 220350
rect 471622 220294 471678 220350
rect 471250 220170 471306 220226
rect 471374 220170 471430 220226
rect 471498 220170 471554 220226
rect 471622 220170 471678 220226
rect 471250 220046 471306 220102
rect 471374 220046 471430 220102
rect 471498 220046 471554 220102
rect 471622 220046 471678 220102
rect 471250 219922 471306 219978
rect 471374 219922 471430 219978
rect 471498 219922 471554 219978
rect 471622 219922 471678 219978
rect 471250 202294 471306 202350
rect 471374 202294 471430 202350
rect 471498 202294 471554 202350
rect 471622 202294 471678 202350
rect 471250 202170 471306 202226
rect 471374 202170 471430 202226
rect 471498 202170 471554 202226
rect 471622 202170 471678 202226
rect 471250 202046 471306 202102
rect 471374 202046 471430 202102
rect 471498 202046 471554 202102
rect 471622 202046 471678 202102
rect 471250 201922 471306 201978
rect 471374 201922 471430 201978
rect 471498 201922 471554 201978
rect 471622 201922 471678 201978
rect 471250 184294 471306 184350
rect 471374 184294 471430 184350
rect 471498 184294 471554 184350
rect 471622 184294 471678 184350
rect 471250 184170 471306 184226
rect 471374 184170 471430 184226
rect 471498 184170 471554 184226
rect 471622 184170 471678 184226
rect 471250 184046 471306 184102
rect 471374 184046 471430 184102
rect 471498 184046 471554 184102
rect 471622 184046 471678 184102
rect 471250 183922 471306 183978
rect 471374 183922 471430 183978
rect 471498 183922 471554 183978
rect 471622 183922 471678 183978
rect 471250 166294 471306 166350
rect 471374 166294 471430 166350
rect 471498 166294 471554 166350
rect 471622 166294 471678 166350
rect 471250 166170 471306 166226
rect 471374 166170 471430 166226
rect 471498 166170 471554 166226
rect 471622 166170 471678 166226
rect 471250 166046 471306 166102
rect 471374 166046 471430 166102
rect 471498 166046 471554 166102
rect 471622 166046 471678 166102
rect 471250 165922 471306 165978
rect 471374 165922 471430 165978
rect 471498 165922 471554 165978
rect 471622 165922 471678 165978
rect 471250 148294 471306 148350
rect 471374 148294 471430 148350
rect 471498 148294 471554 148350
rect 471622 148294 471678 148350
rect 471250 148170 471306 148226
rect 471374 148170 471430 148226
rect 471498 148170 471554 148226
rect 471622 148170 471678 148226
rect 471250 148046 471306 148102
rect 471374 148046 471430 148102
rect 471498 148046 471554 148102
rect 471622 148046 471678 148102
rect 471250 147922 471306 147978
rect 471374 147922 471430 147978
rect 471498 147922 471554 147978
rect 471622 147922 471678 147978
rect 471250 130294 471306 130350
rect 471374 130294 471430 130350
rect 471498 130294 471554 130350
rect 471622 130294 471678 130350
rect 471250 130170 471306 130226
rect 471374 130170 471430 130226
rect 471498 130170 471554 130226
rect 471622 130170 471678 130226
rect 471250 130046 471306 130102
rect 471374 130046 471430 130102
rect 471498 130046 471554 130102
rect 471622 130046 471678 130102
rect 471250 129922 471306 129978
rect 471374 129922 471430 129978
rect 471498 129922 471554 129978
rect 471622 129922 471678 129978
rect 471250 112294 471306 112350
rect 471374 112294 471430 112350
rect 471498 112294 471554 112350
rect 471622 112294 471678 112350
rect 471250 112170 471306 112226
rect 471374 112170 471430 112226
rect 471498 112170 471554 112226
rect 471622 112170 471678 112226
rect 471250 112046 471306 112102
rect 471374 112046 471430 112102
rect 471498 112046 471554 112102
rect 471622 112046 471678 112102
rect 471250 111922 471306 111978
rect 471374 111922 471430 111978
rect 471498 111922 471554 111978
rect 471622 111922 471678 111978
rect 471250 94294 471306 94350
rect 471374 94294 471430 94350
rect 471498 94294 471554 94350
rect 471622 94294 471678 94350
rect 471250 94170 471306 94226
rect 471374 94170 471430 94226
rect 471498 94170 471554 94226
rect 471622 94170 471678 94226
rect 471250 94046 471306 94102
rect 471374 94046 471430 94102
rect 471498 94046 471554 94102
rect 471622 94046 471678 94102
rect 471250 93922 471306 93978
rect 471374 93922 471430 93978
rect 471498 93922 471554 93978
rect 471622 93922 471678 93978
rect 471250 76294 471306 76350
rect 471374 76294 471430 76350
rect 471498 76294 471554 76350
rect 471622 76294 471678 76350
rect 471250 76170 471306 76226
rect 471374 76170 471430 76226
rect 471498 76170 471554 76226
rect 471622 76170 471678 76226
rect 471250 76046 471306 76102
rect 471374 76046 471430 76102
rect 471498 76046 471554 76102
rect 471622 76046 471678 76102
rect 471250 75922 471306 75978
rect 471374 75922 471430 75978
rect 471498 75922 471554 75978
rect 471622 75922 471678 75978
rect 471250 58294 471306 58350
rect 471374 58294 471430 58350
rect 471498 58294 471554 58350
rect 471622 58294 471678 58350
rect 471250 58170 471306 58226
rect 471374 58170 471430 58226
rect 471498 58170 471554 58226
rect 471622 58170 471678 58226
rect 471250 58046 471306 58102
rect 471374 58046 471430 58102
rect 471498 58046 471554 58102
rect 471622 58046 471678 58102
rect 471250 57922 471306 57978
rect 471374 57922 471430 57978
rect 471498 57922 471554 57978
rect 471622 57922 471678 57978
rect 471250 40294 471306 40350
rect 471374 40294 471430 40350
rect 471498 40294 471554 40350
rect 471622 40294 471678 40350
rect 471250 40170 471306 40226
rect 471374 40170 471430 40226
rect 471498 40170 471554 40226
rect 471622 40170 471678 40226
rect 471250 40046 471306 40102
rect 471374 40046 471430 40102
rect 471498 40046 471554 40102
rect 471622 40046 471678 40102
rect 471250 39922 471306 39978
rect 471374 39922 471430 39978
rect 471498 39922 471554 39978
rect 471622 39922 471678 39978
rect 471250 22294 471306 22350
rect 471374 22294 471430 22350
rect 471498 22294 471554 22350
rect 471622 22294 471678 22350
rect 471250 22170 471306 22226
rect 471374 22170 471430 22226
rect 471498 22170 471554 22226
rect 471622 22170 471678 22226
rect 471250 22046 471306 22102
rect 471374 22046 471430 22102
rect 471498 22046 471554 22102
rect 471622 22046 471678 22102
rect 471250 21922 471306 21978
rect 471374 21922 471430 21978
rect 471498 21922 471554 21978
rect 471622 21922 471678 21978
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 474970 598116 475026 598172
rect 475094 598116 475150 598172
rect 475218 598116 475274 598172
rect 475342 598116 475398 598172
rect 474970 597992 475026 598048
rect 475094 597992 475150 598048
rect 475218 597992 475274 598048
rect 475342 597992 475398 598048
rect 474970 597868 475026 597924
rect 475094 597868 475150 597924
rect 475218 597868 475274 597924
rect 475342 597868 475398 597924
rect 474970 597744 475026 597800
rect 475094 597744 475150 597800
rect 475218 597744 475274 597800
rect 475342 597744 475398 597800
rect 474970 586294 475026 586350
rect 475094 586294 475150 586350
rect 475218 586294 475274 586350
rect 475342 586294 475398 586350
rect 474970 586170 475026 586226
rect 475094 586170 475150 586226
rect 475218 586170 475274 586226
rect 475342 586170 475398 586226
rect 474970 586046 475026 586102
rect 475094 586046 475150 586102
rect 475218 586046 475274 586102
rect 475342 586046 475398 586102
rect 474970 585922 475026 585978
rect 475094 585922 475150 585978
rect 475218 585922 475274 585978
rect 475342 585922 475398 585978
rect 474970 568294 475026 568350
rect 475094 568294 475150 568350
rect 475218 568294 475274 568350
rect 475342 568294 475398 568350
rect 474970 568170 475026 568226
rect 475094 568170 475150 568226
rect 475218 568170 475274 568226
rect 475342 568170 475398 568226
rect 474970 568046 475026 568102
rect 475094 568046 475150 568102
rect 475218 568046 475274 568102
rect 475342 568046 475398 568102
rect 474970 567922 475026 567978
rect 475094 567922 475150 567978
rect 475218 567922 475274 567978
rect 475342 567922 475398 567978
rect 474970 550294 475026 550350
rect 475094 550294 475150 550350
rect 475218 550294 475274 550350
rect 475342 550294 475398 550350
rect 474970 550170 475026 550226
rect 475094 550170 475150 550226
rect 475218 550170 475274 550226
rect 475342 550170 475398 550226
rect 474970 550046 475026 550102
rect 475094 550046 475150 550102
rect 475218 550046 475274 550102
rect 475342 550046 475398 550102
rect 474970 549922 475026 549978
rect 475094 549922 475150 549978
rect 475218 549922 475274 549978
rect 475342 549922 475398 549978
rect 474970 532294 475026 532350
rect 475094 532294 475150 532350
rect 475218 532294 475274 532350
rect 475342 532294 475398 532350
rect 474970 532170 475026 532226
rect 475094 532170 475150 532226
rect 475218 532170 475274 532226
rect 475342 532170 475398 532226
rect 474970 532046 475026 532102
rect 475094 532046 475150 532102
rect 475218 532046 475274 532102
rect 475342 532046 475398 532102
rect 474970 531922 475026 531978
rect 475094 531922 475150 531978
rect 475218 531922 475274 531978
rect 475342 531922 475398 531978
rect 474970 514294 475026 514350
rect 475094 514294 475150 514350
rect 475218 514294 475274 514350
rect 475342 514294 475398 514350
rect 474970 514170 475026 514226
rect 475094 514170 475150 514226
rect 475218 514170 475274 514226
rect 475342 514170 475398 514226
rect 474970 514046 475026 514102
rect 475094 514046 475150 514102
rect 475218 514046 475274 514102
rect 475342 514046 475398 514102
rect 474970 513922 475026 513978
rect 475094 513922 475150 513978
rect 475218 513922 475274 513978
rect 475342 513922 475398 513978
rect 474970 496294 475026 496350
rect 475094 496294 475150 496350
rect 475218 496294 475274 496350
rect 475342 496294 475398 496350
rect 474970 496170 475026 496226
rect 475094 496170 475150 496226
rect 475218 496170 475274 496226
rect 475342 496170 475398 496226
rect 474970 496046 475026 496102
rect 475094 496046 475150 496102
rect 475218 496046 475274 496102
rect 475342 496046 475398 496102
rect 474970 495922 475026 495978
rect 475094 495922 475150 495978
rect 475218 495922 475274 495978
rect 475342 495922 475398 495978
rect 474970 478294 475026 478350
rect 475094 478294 475150 478350
rect 475218 478294 475274 478350
rect 475342 478294 475398 478350
rect 474970 478170 475026 478226
rect 475094 478170 475150 478226
rect 475218 478170 475274 478226
rect 475342 478170 475398 478226
rect 474970 478046 475026 478102
rect 475094 478046 475150 478102
rect 475218 478046 475274 478102
rect 475342 478046 475398 478102
rect 474970 477922 475026 477978
rect 475094 477922 475150 477978
rect 475218 477922 475274 477978
rect 475342 477922 475398 477978
rect 474970 460294 475026 460350
rect 475094 460294 475150 460350
rect 475218 460294 475274 460350
rect 475342 460294 475398 460350
rect 474970 460170 475026 460226
rect 475094 460170 475150 460226
rect 475218 460170 475274 460226
rect 475342 460170 475398 460226
rect 474970 460046 475026 460102
rect 475094 460046 475150 460102
rect 475218 460046 475274 460102
rect 475342 460046 475398 460102
rect 474970 459922 475026 459978
rect 475094 459922 475150 459978
rect 475218 459922 475274 459978
rect 475342 459922 475398 459978
rect 474970 442294 475026 442350
rect 475094 442294 475150 442350
rect 475218 442294 475274 442350
rect 475342 442294 475398 442350
rect 474970 442170 475026 442226
rect 475094 442170 475150 442226
rect 475218 442170 475274 442226
rect 475342 442170 475398 442226
rect 474970 442046 475026 442102
rect 475094 442046 475150 442102
rect 475218 442046 475274 442102
rect 475342 442046 475398 442102
rect 474970 441922 475026 441978
rect 475094 441922 475150 441978
rect 475218 441922 475274 441978
rect 475342 441922 475398 441978
rect 474970 424294 475026 424350
rect 475094 424294 475150 424350
rect 475218 424294 475274 424350
rect 475342 424294 475398 424350
rect 474970 424170 475026 424226
rect 475094 424170 475150 424226
rect 475218 424170 475274 424226
rect 475342 424170 475398 424226
rect 474970 424046 475026 424102
rect 475094 424046 475150 424102
rect 475218 424046 475274 424102
rect 475342 424046 475398 424102
rect 474970 423922 475026 423978
rect 475094 423922 475150 423978
rect 475218 423922 475274 423978
rect 475342 423922 475398 423978
rect 474970 406294 475026 406350
rect 475094 406294 475150 406350
rect 475218 406294 475274 406350
rect 475342 406294 475398 406350
rect 474970 406170 475026 406226
rect 475094 406170 475150 406226
rect 475218 406170 475274 406226
rect 475342 406170 475398 406226
rect 474970 406046 475026 406102
rect 475094 406046 475150 406102
rect 475218 406046 475274 406102
rect 475342 406046 475398 406102
rect 474970 405922 475026 405978
rect 475094 405922 475150 405978
rect 475218 405922 475274 405978
rect 475342 405922 475398 405978
rect 474970 388294 475026 388350
rect 475094 388294 475150 388350
rect 475218 388294 475274 388350
rect 475342 388294 475398 388350
rect 474970 388170 475026 388226
rect 475094 388170 475150 388226
rect 475218 388170 475274 388226
rect 475342 388170 475398 388226
rect 474970 388046 475026 388102
rect 475094 388046 475150 388102
rect 475218 388046 475274 388102
rect 475342 388046 475398 388102
rect 474970 387922 475026 387978
rect 475094 387922 475150 387978
rect 475218 387922 475274 387978
rect 475342 387922 475398 387978
rect 474970 370294 475026 370350
rect 475094 370294 475150 370350
rect 475218 370294 475274 370350
rect 475342 370294 475398 370350
rect 474970 370170 475026 370226
rect 475094 370170 475150 370226
rect 475218 370170 475274 370226
rect 475342 370170 475398 370226
rect 474970 370046 475026 370102
rect 475094 370046 475150 370102
rect 475218 370046 475274 370102
rect 475342 370046 475398 370102
rect 474970 369922 475026 369978
rect 475094 369922 475150 369978
rect 475218 369922 475274 369978
rect 475342 369922 475398 369978
rect 474970 352294 475026 352350
rect 475094 352294 475150 352350
rect 475218 352294 475274 352350
rect 475342 352294 475398 352350
rect 474970 352170 475026 352226
rect 475094 352170 475150 352226
rect 475218 352170 475274 352226
rect 475342 352170 475398 352226
rect 474970 352046 475026 352102
rect 475094 352046 475150 352102
rect 475218 352046 475274 352102
rect 475342 352046 475398 352102
rect 474970 351922 475026 351978
rect 475094 351922 475150 351978
rect 475218 351922 475274 351978
rect 475342 351922 475398 351978
rect 474970 334294 475026 334350
rect 475094 334294 475150 334350
rect 475218 334294 475274 334350
rect 475342 334294 475398 334350
rect 474970 334170 475026 334226
rect 475094 334170 475150 334226
rect 475218 334170 475274 334226
rect 475342 334170 475398 334226
rect 474970 334046 475026 334102
rect 475094 334046 475150 334102
rect 475218 334046 475274 334102
rect 475342 334046 475398 334102
rect 474970 333922 475026 333978
rect 475094 333922 475150 333978
rect 475218 333922 475274 333978
rect 475342 333922 475398 333978
rect 474970 316294 475026 316350
rect 475094 316294 475150 316350
rect 475218 316294 475274 316350
rect 475342 316294 475398 316350
rect 474970 316170 475026 316226
rect 475094 316170 475150 316226
rect 475218 316170 475274 316226
rect 475342 316170 475398 316226
rect 474970 316046 475026 316102
rect 475094 316046 475150 316102
rect 475218 316046 475274 316102
rect 475342 316046 475398 316102
rect 474970 315922 475026 315978
rect 475094 315922 475150 315978
rect 475218 315922 475274 315978
rect 475342 315922 475398 315978
rect 474970 298294 475026 298350
rect 475094 298294 475150 298350
rect 475218 298294 475274 298350
rect 475342 298294 475398 298350
rect 474970 298170 475026 298226
rect 475094 298170 475150 298226
rect 475218 298170 475274 298226
rect 475342 298170 475398 298226
rect 474970 298046 475026 298102
rect 475094 298046 475150 298102
rect 475218 298046 475274 298102
rect 475342 298046 475398 298102
rect 474970 297922 475026 297978
rect 475094 297922 475150 297978
rect 475218 297922 475274 297978
rect 475342 297922 475398 297978
rect 474970 280294 475026 280350
rect 475094 280294 475150 280350
rect 475218 280294 475274 280350
rect 475342 280294 475398 280350
rect 474970 280170 475026 280226
rect 475094 280170 475150 280226
rect 475218 280170 475274 280226
rect 475342 280170 475398 280226
rect 474970 280046 475026 280102
rect 475094 280046 475150 280102
rect 475218 280046 475274 280102
rect 475342 280046 475398 280102
rect 474970 279922 475026 279978
rect 475094 279922 475150 279978
rect 475218 279922 475274 279978
rect 475342 279922 475398 279978
rect 474970 262294 475026 262350
rect 475094 262294 475150 262350
rect 475218 262294 475274 262350
rect 475342 262294 475398 262350
rect 474970 262170 475026 262226
rect 475094 262170 475150 262226
rect 475218 262170 475274 262226
rect 475342 262170 475398 262226
rect 474970 262046 475026 262102
rect 475094 262046 475150 262102
rect 475218 262046 475274 262102
rect 475342 262046 475398 262102
rect 474970 261922 475026 261978
rect 475094 261922 475150 261978
rect 475218 261922 475274 261978
rect 475342 261922 475398 261978
rect 474970 244294 475026 244350
rect 475094 244294 475150 244350
rect 475218 244294 475274 244350
rect 475342 244294 475398 244350
rect 474970 244170 475026 244226
rect 475094 244170 475150 244226
rect 475218 244170 475274 244226
rect 475342 244170 475398 244226
rect 474970 244046 475026 244102
rect 475094 244046 475150 244102
rect 475218 244046 475274 244102
rect 475342 244046 475398 244102
rect 474970 243922 475026 243978
rect 475094 243922 475150 243978
rect 475218 243922 475274 243978
rect 475342 243922 475398 243978
rect 474970 226294 475026 226350
rect 475094 226294 475150 226350
rect 475218 226294 475274 226350
rect 475342 226294 475398 226350
rect 474970 226170 475026 226226
rect 475094 226170 475150 226226
rect 475218 226170 475274 226226
rect 475342 226170 475398 226226
rect 474970 226046 475026 226102
rect 475094 226046 475150 226102
rect 475218 226046 475274 226102
rect 475342 226046 475398 226102
rect 474970 225922 475026 225978
rect 475094 225922 475150 225978
rect 475218 225922 475274 225978
rect 475342 225922 475398 225978
rect 474970 208294 475026 208350
rect 475094 208294 475150 208350
rect 475218 208294 475274 208350
rect 475342 208294 475398 208350
rect 474970 208170 475026 208226
rect 475094 208170 475150 208226
rect 475218 208170 475274 208226
rect 475342 208170 475398 208226
rect 474970 208046 475026 208102
rect 475094 208046 475150 208102
rect 475218 208046 475274 208102
rect 475342 208046 475398 208102
rect 474970 207922 475026 207978
rect 475094 207922 475150 207978
rect 475218 207922 475274 207978
rect 475342 207922 475398 207978
rect 474970 190294 475026 190350
rect 475094 190294 475150 190350
rect 475218 190294 475274 190350
rect 475342 190294 475398 190350
rect 474970 190170 475026 190226
rect 475094 190170 475150 190226
rect 475218 190170 475274 190226
rect 475342 190170 475398 190226
rect 474970 190046 475026 190102
rect 475094 190046 475150 190102
rect 475218 190046 475274 190102
rect 475342 190046 475398 190102
rect 474970 189922 475026 189978
rect 475094 189922 475150 189978
rect 475218 189922 475274 189978
rect 475342 189922 475398 189978
rect 474970 172294 475026 172350
rect 475094 172294 475150 172350
rect 475218 172294 475274 172350
rect 475342 172294 475398 172350
rect 474970 172170 475026 172226
rect 475094 172170 475150 172226
rect 475218 172170 475274 172226
rect 475342 172170 475398 172226
rect 474970 172046 475026 172102
rect 475094 172046 475150 172102
rect 475218 172046 475274 172102
rect 475342 172046 475398 172102
rect 474970 171922 475026 171978
rect 475094 171922 475150 171978
rect 475218 171922 475274 171978
rect 475342 171922 475398 171978
rect 474970 154294 475026 154350
rect 475094 154294 475150 154350
rect 475218 154294 475274 154350
rect 475342 154294 475398 154350
rect 474970 154170 475026 154226
rect 475094 154170 475150 154226
rect 475218 154170 475274 154226
rect 475342 154170 475398 154226
rect 474970 154046 475026 154102
rect 475094 154046 475150 154102
rect 475218 154046 475274 154102
rect 475342 154046 475398 154102
rect 474970 153922 475026 153978
rect 475094 153922 475150 153978
rect 475218 153922 475274 153978
rect 475342 153922 475398 153978
rect 474970 136294 475026 136350
rect 475094 136294 475150 136350
rect 475218 136294 475274 136350
rect 475342 136294 475398 136350
rect 474970 136170 475026 136226
rect 475094 136170 475150 136226
rect 475218 136170 475274 136226
rect 475342 136170 475398 136226
rect 474970 136046 475026 136102
rect 475094 136046 475150 136102
rect 475218 136046 475274 136102
rect 475342 136046 475398 136102
rect 474970 135922 475026 135978
rect 475094 135922 475150 135978
rect 475218 135922 475274 135978
rect 475342 135922 475398 135978
rect 474970 118294 475026 118350
rect 475094 118294 475150 118350
rect 475218 118294 475274 118350
rect 475342 118294 475398 118350
rect 474970 118170 475026 118226
rect 475094 118170 475150 118226
rect 475218 118170 475274 118226
rect 475342 118170 475398 118226
rect 474970 118046 475026 118102
rect 475094 118046 475150 118102
rect 475218 118046 475274 118102
rect 475342 118046 475398 118102
rect 474970 117922 475026 117978
rect 475094 117922 475150 117978
rect 475218 117922 475274 117978
rect 475342 117922 475398 117978
rect 474970 100294 475026 100350
rect 475094 100294 475150 100350
rect 475218 100294 475274 100350
rect 475342 100294 475398 100350
rect 474970 100170 475026 100226
rect 475094 100170 475150 100226
rect 475218 100170 475274 100226
rect 475342 100170 475398 100226
rect 474970 100046 475026 100102
rect 475094 100046 475150 100102
rect 475218 100046 475274 100102
rect 475342 100046 475398 100102
rect 474970 99922 475026 99978
rect 475094 99922 475150 99978
rect 475218 99922 475274 99978
rect 475342 99922 475398 99978
rect 474970 82294 475026 82350
rect 475094 82294 475150 82350
rect 475218 82294 475274 82350
rect 475342 82294 475398 82350
rect 474970 82170 475026 82226
rect 475094 82170 475150 82226
rect 475218 82170 475274 82226
rect 475342 82170 475398 82226
rect 474970 82046 475026 82102
rect 475094 82046 475150 82102
rect 475218 82046 475274 82102
rect 475342 82046 475398 82102
rect 474970 81922 475026 81978
rect 475094 81922 475150 81978
rect 475218 81922 475274 81978
rect 475342 81922 475398 81978
rect 474970 64294 475026 64350
rect 475094 64294 475150 64350
rect 475218 64294 475274 64350
rect 475342 64294 475398 64350
rect 474970 64170 475026 64226
rect 475094 64170 475150 64226
rect 475218 64170 475274 64226
rect 475342 64170 475398 64226
rect 474970 64046 475026 64102
rect 475094 64046 475150 64102
rect 475218 64046 475274 64102
rect 475342 64046 475398 64102
rect 474970 63922 475026 63978
rect 475094 63922 475150 63978
rect 475218 63922 475274 63978
rect 475342 63922 475398 63978
rect 474970 46294 475026 46350
rect 475094 46294 475150 46350
rect 475218 46294 475274 46350
rect 475342 46294 475398 46350
rect 474970 46170 475026 46226
rect 475094 46170 475150 46226
rect 475218 46170 475274 46226
rect 475342 46170 475398 46226
rect 474970 46046 475026 46102
rect 475094 46046 475150 46102
rect 475218 46046 475274 46102
rect 475342 46046 475398 46102
rect 474970 45922 475026 45978
rect 475094 45922 475150 45978
rect 475218 45922 475274 45978
rect 475342 45922 475398 45978
rect 474970 28294 475026 28350
rect 475094 28294 475150 28350
rect 475218 28294 475274 28350
rect 475342 28294 475398 28350
rect 474970 28170 475026 28226
rect 475094 28170 475150 28226
rect 475218 28170 475274 28226
rect 475342 28170 475398 28226
rect 474970 28046 475026 28102
rect 475094 28046 475150 28102
rect 475218 28046 475274 28102
rect 475342 28046 475398 28102
rect 474970 27922 475026 27978
rect 475094 27922 475150 27978
rect 475218 27922 475274 27978
rect 475342 27922 475398 27978
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 489250 526294 489306 526350
rect 489374 526294 489430 526350
rect 489498 526294 489554 526350
rect 489622 526294 489678 526350
rect 489250 526170 489306 526226
rect 489374 526170 489430 526226
rect 489498 526170 489554 526226
rect 489622 526170 489678 526226
rect 489250 526046 489306 526102
rect 489374 526046 489430 526102
rect 489498 526046 489554 526102
rect 489622 526046 489678 526102
rect 489250 525922 489306 525978
rect 489374 525922 489430 525978
rect 489498 525922 489554 525978
rect 489622 525922 489678 525978
rect 489250 508294 489306 508350
rect 489374 508294 489430 508350
rect 489498 508294 489554 508350
rect 489622 508294 489678 508350
rect 489250 508170 489306 508226
rect 489374 508170 489430 508226
rect 489498 508170 489554 508226
rect 489622 508170 489678 508226
rect 489250 508046 489306 508102
rect 489374 508046 489430 508102
rect 489498 508046 489554 508102
rect 489622 508046 489678 508102
rect 489250 507922 489306 507978
rect 489374 507922 489430 507978
rect 489498 507922 489554 507978
rect 489622 507922 489678 507978
rect 489250 490294 489306 490350
rect 489374 490294 489430 490350
rect 489498 490294 489554 490350
rect 489622 490294 489678 490350
rect 489250 490170 489306 490226
rect 489374 490170 489430 490226
rect 489498 490170 489554 490226
rect 489622 490170 489678 490226
rect 489250 490046 489306 490102
rect 489374 490046 489430 490102
rect 489498 490046 489554 490102
rect 489622 490046 489678 490102
rect 489250 489922 489306 489978
rect 489374 489922 489430 489978
rect 489498 489922 489554 489978
rect 489622 489922 489678 489978
rect 489250 472294 489306 472350
rect 489374 472294 489430 472350
rect 489498 472294 489554 472350
rect 489622 472294 489678 472350
rect 489250 472170 489306 472226
rect 489374 472170 489430 472226
rect 489498 472170 489554 472226
rect 489622 472170 489678 472226
rect 489250 472046 489306 472102
rect 489374 472046 489430 472102
rect 489498 472046 489554 472102
rect 489622 472046 489678 472102
rect 489250 471922 489306 471978
rect 489374 471922 489430 471978
rect 489498 471922 489554 471978
rect 489622 471922 489678 471978
rect 489250 454294 489306 454350
rect 489374 454294 489430 454350
rect 489498 454294 489554 454350
rect 489622 454294 489678 454350
rect 489250 454170 489306 454226
rect 489374 454170 489430 454226
rect 489498 454170 489554 454226
rect 489622 454170 489678 454226
rect 489250 454046 489306 454102
rect 489374 454046 489430 454102
rect 489498 454046 489554 454102
rect 489622 454046 489678 454102
rect 489250 453922 489306 453978
rect 489374 453922 489430 453978
rect 489498 453922 489554 453978
rect 489622 453922 489678 453978
rect 489250 436294 489306 436350
rect 489374 436294 489430 436350
rect 489498 436294 489554 436350
rect 489622 436294 489678 436350
rect 489250 436170 489306 436226
rect 489374 436170 489430 436226
rect 489498 436170 489554 436226
rect 489622 436170 489678 436226
rect 489250 436046 489306 436102
rect 489374 436046 489430 436102
rect 489498 436046 489554 436102
rect 489622 436046 489678 436102
rect 489250 435922 489306 435978
rect 489374 435922 489430 435978
rect 489498 435922 489554 435978
rect 489622 435922 489678 435978
rect 489250 418294 489306 418350
rect 489374 418294 489430 418350
rect 489498 418294 489554 418350
rect 489622 418294 489678 418350
rect 489250 418170 489306 418226
rect 489374 418170 489430 418226
rect 489498 418170 489554 418226
rect 489622 418170 489678 418226
rect 489250 418046 489306 418102
rect 489374 418046 489430 418102
rect 489498 418046 489554 418102
rect 489622 418046 489678 418102
rect 489250 417922 489306 417978
rect 489374 417922 489430 417978
rect 489498 417922 489554 417978
rect 489622 417922 489678 417978
rect 489250 400294 489306 400350
rect 489374 400294 489430 400350
rect 489498 400294 489554 400350
rect 489622 400294 489678 400350
rect 489250 400170 489306 400226
rect 489374 400170 489430 400226
rect 489498 400170 489554 400226
rect 489622 400170 489678 400226
rect 489250 400046 489306 400102
rect 489374 400046 489430 400102
rect 489498 400046 489554 400102
rect 489622 400046 489678 400102
rect 489250 399922 489306 399978
rect 489374 399922 489430 399978
rect 489498 399922 489554 399978
rect 489622 399922 489678 399978
rect 489250 382294 489306 382350
rect 489374 382294 489430 382350
rect 489498 382294 489554 382350
rect 489622 382294 489678 382350
rect 489250 382170 489306 382226
rect 489374 382170 489430 382226
rect 489498 382170 489554 382226
rect 489622 382170 489678 382226
rect 489250 382046 489306 382102
rect 489374 382046 489430 382102
rect 489498 382046 489554 382102
rect 489622 382046 489678 382102
rect 489250 381922 489306 381978
rect 489374 381922 489430 381978
rect 489498 381922 489554 381978
rect 489622 381922 489678 381978
rect 489250 364294 489306 364350
rect 489374 364294 489430 364350
rect 489498 364294 489554 364350
rect 489622 364294 489678 364350
rect 489250 364170 489306 364226
rect 489374 364170 489430 364226
rect 489498 364170 489554 364226
rect 489622 364170 489678 364226
rect 489250 364046 489306 364102
rect 489374 364046 489430 364102
rect 489498 364046 489554 364102
rect 489622 364046 489678 364102
rect 489250 363922 489306 363978
rect 489374 363922 489430 363978
rect 489498 363922 489554 363978
rect 489622 363922 489678 363978
rect 489250 346294 489306 346350
rect 489374 346294 489430 346350
rect 489498 346294 489554 346350
rect 489622 346294 489678 346350
rect 489250 346170 489306 346226
rect 489374 346170 489430 346226
rect 489498 346170 489554 346226
rect 489622 346170 489678 346226
rect 489250 346046 489306 346102
rect 489374 346046 489430 346102
rect 489498 346046 489554 346102
rect 489622 346046 489678 346102
rect 489250 345922 489306 345978
rect 489374 345922 489430 345978
rect 489498 345922 489554 345978
rect 489622 345922 489678 345978
rect 489250 328294 489306 328350
rect 489374 328294 489430 328350
rect 489498 328294 489554 328350
rect 489622 328294 489678 328350
rect 489250 328170 489306 328226
rect 489374 328170 489430 328226
rect 489498 328170 489554 328226
rect 489622 328170 489678 328226
rect 489250 328046 489306 328102
rect 489374 328046 489430 328102
rect 489498 328046 489554 328102
rect 489622 328046 489678 328102
rect 489250 327922 489306 327978
rect 489374 327922 489430 327978
rect 489498 327922 489554 327978
rect 489622 327922 489678 327978
rect 489250 310294 489306 310350
rect 489374 310294 489430 310350
rect 489498 310294 489554 310350
rect 489622 310294 489678 310350
rect 489250 310170 489306 310226
rect 489374 310170 489430 310226
rect 489498 310170 489554 310226
rect 489622 310170 489678 310226
rect 489250 310046 489306 310102
rect 489374 310046 489430 310102
rect 489498 310046 489554 310102
rect 489622 310046 489678 310102
rect 489250 309922 489306 309978
rect 489374 309922 489430 309978
rect 489498 309922 489554 309978
rect 489622 309922 489678 309978
rect 489250 292294 489306 292350
rect 489374 292294 489430 292350
rect 489498 292294 489554 292350
rect 489622 292294 489678 292350
rect 489250 292170 489306 292226
rect 489374 292170 489430 292226
rect 489498 292170 489554 292226
rect 489622 292170 489678 292226
rect 489250 292046 489306 292102
rect 489374 292046 489430 292102
rect 489498 292046 489554 292102
rect 489622 292046 489678 292102
rect 489250 291922 489306 291978
rect 489374 291922 489430 291978
rect 489498 291922 489554 291978
rect 489622 291922 489678 291978
rect 489250 274294 489306 274350
rect 489374 274294 489430 274350
rect 489498 274294 489554 274350
rect 489622 274294 489678 274350
rect 489250 274170 489306 274226
rect 489374 274170 489430 274226
rect 489498 274170 489554 274226
rect 489622 274170 489678 274226
rect 489250 274046 489306 274102
rect 489374 274046 489430 274102
rect 489498 274046 489554 274102
rect 489622 274046 489678 274102
rect 489250 273922 489306 273978
rect 489374 273922 489430 273978
rect 489498 273922 489554 273978
rect 489622 273922 489678 273978
rect 489250 256294 489306 256350
rect 489374 256294 489430 256350
rect 489498 256294 489554 256350
rect 489622 256294 489678 256350
rect 489250 256170 489306 256226
rect 489374 256170 489430 256226
rect 489498 256170 489554 256226
rect 489622 256170 489678 256226
rect 489250 256046 489306 256102
rect 489374 256046 489430 256102
rect 489498 256046 489554 256102
rect 489622 256046 489678 256102
rect 489250 255922 489306 255978
rect 489374 255922 489430 255978
rect 489498 255922 489554 255978
rect 489622 255922 489678 255978
rect 489250 238294 489306 238350
rect 489374 238294 489430 238350
rect 489498 238294 489554 238350
rect 489622 238294 489678 238350
rect 489250 238170 489306 238226
rect 489374 238170 489430 238226
rect 489498 238170 489554 238226
rect 489622 238170 489678 238226
rect 489250 238046 489306 238102
rect 489374 238046 489430 238102
rect 489498 238046 489554 238102
rect 489622 238046 489678 238102
rect 489250 237922 489306 237978
rect 489374 237922 489430 237978
rect 489498 237922 489554 237978
rect 489622 237922 489678 237978
rect 489250 220294 489306 220350
rect 489374 220294 489430 220350
rect 489498 220294 489554 220350
rect 489622 220294 489678 220350
rect 489250 220170 489306 220226
rect 489374 220170 489430 220226
rect 489498 220170 489554 220226
rect 489622 220170 489678 220226
rect 489250 220046 489306 220102
rect 489374 220046 489430 220102
rect 489498 220046 489554 220102
rect 489622 220046 489678 220102
rect 489250 219922 489306 219978
rect 489374 219922 489430 219978
rect 489498 219922 489554 219978
rect 489622 219922 489678 219978
rect 489250 202294 489306 202350
rect 489374 202294 489430 202350
rect 489498 202294 489554 202350
rect 489622 202294 489678 202350
rect 489250 202170 489306 202226
rect 489374 202170 489430 202226
rect 489498 202170 489554 202226
rect 489622 202170 489678 202226
rect 489250 202046 489306 202102
rect 489374 202046 489430 202102
rect 489498 202046 489554 202102
rect 489622 202046 489678 202102
rect 489250 201922 489306 201978
rect 489374 201922 489430 201978
rect 489498 201922 489554 201978
rect 489622 201922 489678 201978
rect 489250 184294 489306 184350
rect 489374 184294 489430 184350
rect 489498 184294 489554 184350
rect 489622 184294 489678 184350
rect 489250 184170 489306 184226
rect 489374 184170 489430 184226
rect 489498 184170 489554 184226
rect 489622 184170 489678 184226
rect 489250 184046 489306 184102
rect 489374 184046 489430 184102
rect 489498 184046 489554 184102
rect 489622 184046 489678 184102
rect 489250 183922 489306 183978
rect 489374 183922 489430 183978
rect 489498 183922 489554 183978
rect 489622 183922 489678 183978
rect 489250 166294 489306 166350
rect 489374 166294 489430 166350
rect 489498 166294 489554 166350
rect 489622 166294 489678 166350
rect 489250 166170 489306 166226
rect 489374 166170 489430 166226
rect 489498 166170 489554 166226
rect 489622 166170 489678 166226
rect 489250 166046 489306 166102
rect 489374 166046 489430 166102
rect 489498 166046 489554 166102
rect 489622 166046 489678 166102
rect 489250 165922 489306 165978
rect 489374 165922 489430 165978
rect 489498 165922 489554 165978
rect 489622 165922 489678 165978
rect 489250 148294 489306 148350
rect 489374 148294 489430 148350
rect 489498 148294 489554 148350
rect 489622 148294 489678 148350
rect 489250 148170 489306 148226
rect 489374 148170 489430 148226
rect 489498 148170 489554 148226
rect 489622 148170 489678 148226
rect 489250 148046 489306 148102
rect 489374 148046 489430 148102
rect 489498 148046 489554 148102
rect 489622 148046 489678 148102
rect 489250 147922 489306 147978
rect 489374 147922 489430 147978
rect 489498 147922 489554 147978
rect 489622 147922 489678 147978
rect 489250 130294 489306 130350
rect 489374 130294 489430 130350
rect 489498 130294 489554 130350
rect 489622 130294 489678 130350
rect 489250 130170 489306 130226
rect 489374 130170 489430 130226
rect 489498 130170 489554 130226
rect 489622 130170 489678 130226
rect 489250 130046 489306 130102
rect 489374 130046 489430 130102
rect 489498 130046 489554 130102
rect 489622 130046 489678 130102
rect 489250 129922 489306 129978
rect 489374 129922 489430 129978
rect 489498 129922 489554 129978
rect 489622 129922 489678 129978
rect 489250 112294 489306 112350
rect 489374 112294 489430 112350
rect 489498 112294 489554 112350
rect 489622 112294 489678 112350
rect 489250 112170 489306 112226
rect 489374 112170 489430 112226
rect 489498 112170 489554 112226
rect 489622 112170 489678 112226
rect 489250 112046 489306 112102
rect 489374 112046 489430 112102
rect 489498 112046 489554 112102
rect 489622 112046 489678 112102
rect 489250 111922 489306 111978
rect 489374 111922 489430 111978
rect 489498 111922 489554 111978
rect 489622 111922 489678 111978
rect 489250 94294 489306 94350
rect 489374 94294 489430 94350
rect 489498 94294 489554 94350
rect 489622 94294 489678 94350
rect 489250 94170 489306 94226
rect 489374 94170 489430 94226
rect 489498 94170 489554 94226
rect 489622 94170 489678 94226
rect 489250 94046 489306 94102
rect 489374 94046 489430 94102
rect 489498 94046 489554 94102
rect 489622 94046 489678 94102
rect 489250 93922 489306 93978
rect 489374 93922 489430 93978
rect 489498 93922 489554 93978
rect 489622 93922 489678 93978
rect 489250 76294 489306 76350
rect 489374 76294 489430 76350
rect 489498 76294 489554 76350
rect 489622 76294 489678 76350
rect 489250 76170 489306 76226
rect 489374 76170 489430 76226
rect 489498 76170 489554 76226
rect 489622 76170 489678 76226
rect 489250 76046 489306 76102
rect 489374 76046 489430 76102
rect 489498 76046 489554 76102
rect 489622 76046 489678 76102
rect 489250 75922 489306 75978
rect 489374 75922 489430 75978
rect 489498 75922 489554 75978
rect 489622 75922 489678 75978
rect 489250 58294 489306 58350
rect 489374 58294 489430 58350
rect 489498 58294 489554 58350
rect 489622 58294 489678 58350
rect 489250 58170 489306 58226
rect 489374 58170 489430 58226
rect 489498 58170 489554 58226
rect 489622 58170 489678 58226
rect 489250 58046 489306 58102
rect 489374 58046 489430 58102
rect 489498 58046 489554 58102
rect 489622 58046 489678 58102
rect 489250 57922 489306 57978
rect 489374 57922 489430 57978
rect 489498 57922 489554 57978
rect 489622 57922 489678 57978
rect 489250 40294 489306 40350
rect 489374 40294 489430 40350
rect 489498 40294 489554 40350
rect 489622 40294 489678 40350
rect 489250 40170 489306 40226
rect 489374 40170 489430 40226
rect 489498 40170 489554 40226
rect 489622 40170 489678 40226
rect 489250 40046 489306 40102
rect 489374 40046 489430 40102
rect 489498 40046 489554 40102
rect 489622 40046 489678 40102
rect 489250 39922 489306 39978
rect 489374 39922 489430 39978
rect 489498 39922 489554 39978
rect 489622 39922 489678 39978
rect 489250 22294 489306 22350
rect 489374 22294 489430 22350
rect 489498 22294 489554 22350
rect 489622 22294 489678 22350
rect 489250 22170 489306 22226
rect 489374 22170 489430 22226
rect 489498 22170 489554 22226
rect 489622 22170 489678 22226
rect 489250 22046 489306 22102
rect 489374 22046 489430 22102
rect 489498 22046 489554 22102
rect 489622 22046 489678 22102
rect 489250 21922 489306 21978
rect 489374 21922 489430 21978
rect 489498 21922 489554 21978
rect 489622 21922 489678 21978
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 492970 514294 493026 514350
rect 493094 514294 493150 514350
rect 493218 514294 493274 514350
rect 493342 514294 493398 514350
rect 492970 514170 493026 514226
rect 493094 514170 493150 514226
rect 493218 514170 493274 514226
rect 493342 514170 493398 514226
rect 492970 514046 493026 514102
rect 493094 514046 493150 514102
rect 493218 514046 493274 514102
rect 493342 514046 493398 514102
rect 492970 513922 493026 513978
rect 493094 513922 493150 513978
rect 493218 513922 493274 513978
rect 493342 513922 493398 513978
rect 492970 496294 493026 496350
rect 493094 496294 493150 496350
rect 493218 496294 493274 496350
rect 493342 496294 493398 496350
rect 492970 496170 493026 496226
rect 493094 496170 493150 496226
rect 493218 496170 493274 496226
rect 493342 496170 493398 496226
rect 492970 496046 493026 496102
rect 493094 496046 493150 496102
rect 493218 496046 493274 496102
rect 493342 496046 493398 496102
rect 492970 495922 493026 495978
rect 493094 495922 493150 495978
rect 493218 495922 493274 495978
rect 493342 495922 493398 495978
rect 492970 478294 493026 478350
rect 493094 478294 493150 478350
rect 493218 478294 493274 478350
rect 493342 478294 493398 478350
rect 492970 478170 493026 478226
rect 493094 478170 493150 478226
rect 493218 478170 493274 478226
rect 493342 478170 493398 478226
rect 492970 478046 493026 478102
rect 493094 478046 493150 478102
rect 493218 478046 493274 478102
rect 493342 478046 493398 478102
rect 492970 477922 493026 477978
rect 493094 477922 493150 477978
rect 493218 477922 493274 477978
rect 493342 477922 493398 477978
rect 492970 460294 493026 460350
rect 493094 460294 493150 460350
rect 493218 460294 493274 460350
rect 493342 460294 493398 460350
rect 492970 460170 493026 460226
rect 493094 460170 493150 460226
rect 493218 460170 493274 460226
rect 493342 460170 493398 460226
rect 492970 460046 493026 460102
rect 493094 460046 493150 460102
rect 493218 460046 493274 460102
rect 493342 460046 493398 460102
rect 492970 459922 493026 459978
rect 493094 459922 493150 459978
rect 493218 459922 493274 459978
rect 493342 459922 493398 459978
rect 492970 442294 493026 442350
rect 493094 442294 493150 442350
rect 493218 442294 493274 442350
rect 493342 442294 493398 442350
rect 492970 442170 493026 442226
rect 493094 442170 493150 442226
rect 493218 442170 493274 442226
rect 493342 442170 493398 442226
rect 492970 442046 493026 442102
rect 493094 442046 493150 442102
rect 493218 442046 493274 442102
rect 493342 442046 493398 442102
rect 492970 441922 493026 441978
rect 493094 441922 493150 441978
rect 493218 441922 493274 441978
rect 493342 441922 493398 441978
rect 492970 424294 493026 424350
rect 493094 424294 493150 424350
rect 493218 424294 493274 424350
rect 493342 424294 493398 424350
rect 492970 424170 493026 424226
rect 493094 424170 493150 424226
rect 493218 424170 493274 424226
rect 493342 424170 493398 424226
rect 492970 424046 493026 424102
rect 493094 424046 493150 424102
rect 493218 424046 493274 424102
rect 493342 424046 493398 424102
rect 492970 423922 493026 423978
rect 493094 423922 493150 423978
rect 493218 423922 493274 423978
rect 493342 423922 493398 423978
rect 492970 406294 493026 406350
rect 493094 406294 493150 406350
rect 493218 406294 493274 406350
rect 493342 406294 493398 406350
rect 492970 406170 493026 406226
rect 493094 406170 493150 406226
rect 493218 406170 493274 406226
rect 493342 406170 493398 406226
rect 492970 406046 493026 406102
rect 493094 406046 493150 406102
rect 493218 406046 493274 406102
rect 493342 406046 493398 406102
rect 492970 405922 493026 405978
rect 493094 405922 493150 405978
rect 493218 405922 493274 405978
rect 493342 405922 493398 405978
rect 492970 388294 493026 388350
rect 493094 388294 493150 388350
rect 493218 388294 493274 388350
rect 493342 388294 493398 388350
rect 492970 388170 493026 388226
rect 493094 388170 493150 388226
rect 493218 388170 493274 388226
rect 493342 388170 493398 388226
rect 492970 388046 493026 388102
rect 493094 388046 493150 388102
rect 493218 388046 493274 388102
rect 493342 388046 493398 388102
rect 492970 387922 493026 387978
rect 493094 387922 493150 387978
rect 493218 387922 493274 387978
rect 493342 387922 493398 387978
rect 492970 370294 493026 370350
rect 493094 370294 493150 370350
rect 493218 370294 493274 370350
rect 493342 370294 493398 370350
rect 492970 370170 493026 370226
rect 493094 370170 493150 370226
rect 493218 370170 493274 370226
rect 493342 370170 493398 370226
rect 492970 370046 493026 370102
rect 493094 370046 493150 370102
rect 493218 370046 493274 370102
rect 493342 370046 493398 370102
rect 492970 369922 493026 369978
rect 493094 369922 493150 369978
rect 493218 369922 493274 369978
rect 493342 369922 493398 369978
rect 492970 352294 493026 352350
rect 493094 352294 493150 352350
rect 493218 352294 493274 352350
rect 493342 352294 493398 352350
rect 492970 352170 493026 352226
rect 493094 352170 493150 352226
rect 493218 352170 493274 352226
rect 493342 352170 493398 352226
rect 492970 352046 493026 352102
rect 493094 352046 493150 352102
rect 493218 352046 493274 352102
rect 493342 352046 493398 352102
rect 492970 351922 493026 351978
rect 493094 351922 493150 351978
rect 493218 351922 493274 351978
rect 493342 351922 493398 351978
rect 492970 334294 493026 334350
rect 493094 334294 493150 334350
rect 493218 334294 493274 334350
rect 493342 334294 493398 334350
rect 492970 334170 493026 334226
rect 493094 334170 493150 334226
rect 493218 334170 493274 334226
rect 493342 334170 493398 334226
rect 492970 334046 493026 334102
rect 493094 334046 493150 334102
rect 493218 334046 493274 334102
rect 493342 334046 493398 334102
rect 492970 333922 493026 333978
rect 493094 333922 493150 333978
rect 493218 333922 493274 333978
rect 493342 333922 493398 333978
rect 492970 316294 493026 316350
rect 493094 316294 493150 316350
rect 493218 316294 493274 316350
rect 493342 316294 493398 316350
rect 492970 316170 493026 316226
rect 493094 316170 493150 316226
rect 493218 316170 493274 316226
rect 493342 316170 493398 316226
rect 492970 316046 493026 316102
rect 493094 316046 493150 316102
rect 493218 316046 493274 316102
rect 493342 316046 493398 316102
rect 492970 315922 493026 315978
rect 493094 315922 493150 315978
rect 493218 315922 493274 315978
rect 493342 315922 493398 315978
rect 492970 298294 493026 298350
rect 493094 298294 493150 298350
rect 493218 298294 493274 298350
rect 493342 298294 493398 298350
rect 492970 298170 493026 298226
rect 493094 298170 493150 298226
rect 493218 298170 493274 298226
rect 493342 298170 493398 298226
rect 492970 298046 493026 298102
rect 493094 298046 493150 298102
rect 493218 298046 493274 298102
rect 493342 298046 493398 298102
rect 492970 297922 493026 297978
rect 493094 297922 493150 297978
rect 493218 297922 493274 297978
rect 493342 297922 493398 297978
rect 492970 280294 493026 280350
rect 493094 280294 493150 280350
rect 493218 280294 493274 280350
rect 493342 280294 493398 280350
rect 492970 280170 493026 280226
rect 493094 280170 493150 280226
rect 493218 280170 493274 280226
rect 493342 280170 493398 280226
rect 492970 280046 493026 280102
rect 493094 280046 493150 280102
rect 493218 280046 493274 280102
rect 493342 280046 493398 280102
rect 492970 279922 493026 279978
rect 493094 279922 493150 279978
rect 493218 279922 493274 279978
rect 493342 279922 493398 279978
rect 492970 262294 493026 262350
rect 493094 262294 493150 262350
rect 493218 262294 493274 262350
rect 493342 262294 493398 262350
rect 492970 262170 493026 262226
rect 493094 262170 493150 262226
rect 493218 262170 493274 262226
rect 493342 262170 493398 262226
rect 492970 262046 493026 262102
rect 493094 262046 493150 262102
rect 493218 262046 493274 262102
rect 493342 262046 493398 262102
rect 492970 261922 493026 261978
rect 493094 261922 493150 261978
rect 493218 261922 493274 261978
rect 493342 261922 493398 261978
rect 492970 244294 493026 244350
rect 493094 244294 493150 244350
rect 493218 244294 493274 244350
rect 493342 244294 493398 244350
rect 492970 244170 493026 244226
rect 493094 244170 493150 244226
rect 493218 244170 493274 244226
rect 493342 244170 493398 244226
rect 492970 244046 493026 244102
rect 493094 244046 493150 244102
rect 493218 244046 493274 244102
rect 493342 244046 493398 244102
rect 492970 243922 493026 243978
rect 493094 243922 493150 243978
rect 493218 243922 493274 243978
rect 493342 243922 493398 243978
rect 492970 226294 493026 226350
rect 493094 226294 493150 226350
rect 493218 226294 493274 226350
rect 493342 226294 493398 226350
rect 492970 226170 493026 226226
rect 493094 226170 493150 226226
rect 493218 226170 493274 226226
rect 493342 226170 493398 226226
rect 492970 226046 493026 226102
rect 493094 226046 493150 226102
rect 493218 226046 493274 226102
rect 493342 226046 493398 226102
rect 492970 225922 493026 225978
rect 493094 225922 493150 225978
rect 493218 225922 493274 225978
rect 493342 225922 493398 225978
rect 492970 208294 493026 208350
rect 493094 208294 493150 208350
rect 493218 208294 493274 208350
rect 493342 208294 493398 208350
rect 492970 208170 493026 208226
rect 493094 208170 493150 208226
rect 493218 208170 493274 208226
rect 493342 208170 493398 208226
rect 492970 208046 493026 208102
rect 493094 208046 493150 208102
rect 493218 208046 493274 208102
rect 493342 208046 493398 208102
rect 492970 207922 493026 207978
rect 493094 207922 493150 207978
rect 493218 207922 493274 207978
rect 493342 207922 493398 207978
rect 492970 190294 493026 190350
rect 493094 190294 493150 190350
rect 493218 190294 493274 190350
rect 493342 190294 493398 190350
rect 492970 190170 493026 190226
rect 493094 190170 493150 190226
rect 493218 190170 493274 190226
rect 493342 190170 493398 190226
rect 492970 190046 493026 190102
rect 493094 190046 493150 190102
rect 493218 190046 493274 190102
rect 493342 190046 493398 190102
rect 492970 189922 493026 189978
rect 493094 189922 493150 189978
rect 493218 189922 493274 189978
rect 493342 189922 493398 189978
rect 492970 172294 493026 172350
rect 493094 172294 493150 172350
rect 493218 172294 493274 172350
rect 493342 172294 493398 172350
rect 492970 172170 493026 172226
rect 493094 172170 493150 172226
rect 493218 172170 493274 172226
rect 493342 172170 493398 172226
rect 492970 172046 493026 172102
rect 493094 172046 493150 172102
rect 493218 172046 493274 172102
rect 493342 172046 493398 172102
rect 492970 171922 493026 171978
rect 493094 171922 493150 171978
rect 493218 171922 493274 171978
rect 493342 171922 493398 171978
rect 492970 154294 493026 154350
rect 493094 154294 493150 154350
rect 493218 154294 493274 154350
rect 493342 154294 493398 154350
rect 492970 154170 493026 154226
rect 493094 154170 493150 154226
rect 493218 154170 493274 154226
rect 493342 154170 493398 154226
rect 492970 154046 493026 154102
rect 493094 154046 493150 154102
rect 493218 154046 493274 154102
rect 493342 154046 493398 154102
rect 492970 153922 493026 153978
rect 493094 153922 493150 153978
rect 493218 153922 493274 153978
rect 493342 153922 493398 153978
rect 492970 136294 493026 136350
rect 493094 136294 493150 136350
rect 493218 136294 493274 136350
rect 493342 136294 493398 136350
rect 492970 136170 493026 136226
rect 493094 136170 493150 136226
rect 493218 136170 493274 136226
rect 493342 136170 493398 136226
rect 492970 136046 493026 136102
rect 493094 136046 493150 136102
rect 493218 136046 493274 136102
rect 493342 136046 493398 136102
rect 492970 135922 493026 135978
rect 493094 135922 493150 135978
rect 493218 135922 493274 135978
rect 493342 135922 493398 135978
rect 492970 118294 493026 118350
rect 493094 118294 493150 118350
rect 493218 118294 493274 118350
rect 493342 118294 493398 118350
rect 492970 118170 493026 118226
rect 493094 118170 493150 118226
rect 493218 118170 493274 118226
rect 493342 118170 493398 118226
rect 492970 118046 493026 118102
rect 493094 118046 493150 118102
rect 493218 118046 493274 118102
rect 493342 118046 493398 118102
rect 492970 117922 493026 117978
rect 493094 117922 493150 117978
rect 493218 117922 493274 117978
rect 493342 117922 493398 117978
rect 492970 100294 493026 100350
rect 493094 100294 493150 100350
rect 493218 100294 493274 100350
rect 493342 100294 493398 100350
rect 492970 100170 493026 100226
rect 493094 100170 493150 100226
rect 493218 100170 493274 100226
rect 493342 100170 493398 100226
rect 492970 100046 493026 100102
rect 493094 100046 493150 100102
rect 493218 100046 493274 100102
rect 493342 100046 493398 100102
rect 492970 99922 493026 99978
rect 493094 99922 493150 99978
rect 493218 99922 493274 99978
rect 493342 99922 493398 99978
rect 492970 82294 493026 82350
rect 493094 82294 493150 82350
rect 493218 82294 493274 82350
rect 493342 82294 493398 82350
rect 492970 82170 493026 82226
rect 493094 82170 493150 82226
rect 493218 82170 493274 82226
rect 493342 82170 493398 82226
rect 492970 82046 493026 82102
rect 493094 82046 493150 82102
rect 493218 82046 493274 82102
rect 493342 82046 493398 82102
rect 492970 81922 493026 81978
rect 493094 81922 493150 81978
rect 493218 81922 493274 81978
rect 493342 81922 493398 81978
rect 492970 64294 493026 64350
rect 493094 64294 493150 64350
rect 493218 64294 493274 64350
rect 493342 64294 493398 64350
rect 492970 64170 493026 64226
rect 493094 64170 493150 64226
rect 493218 64170 493274 64226
rect 493342 64170 493398 64226
rect 492970 64046 493026 64102
rect 493094 64046 493150 64102
rect 493218 64046 493274 64102
rect 493342 64046 493398 64102
rect 492970 63922 493026 63978
rect 493094 63922 493150 63978
rect 493218 63922 493274 63978
rect 493342 63922 493398 63978
rect 492970 46294 493026 46350
rect 493094 46294 493150 46350
rect 493218 46294 493274 46350
rect 493342 46294 493398 46350
rect 492970 46170 493026 46226
rect 493094 46170 493150 46226
rect 493218 46170 493274 46226
rect 493342 46170 493398 46226
rect 492970 46046 493026 46102
rect 493094 46046 493150 46102
rect 493218 46046 493274 46102
rect 493342 46046 493398 46102
rect 492970 45922 493026 45978
rect 493094 45922 493150 45978
rect 493218 45922 493274 45978
rect 493342 45922 493398 45978
rect 492970 28294 493026 28350
rect 493094 28294 493150 28350
rect 493218 28294 493274 28350
rect 493342 28294 493398 28350
rect 492970 28170 493026 28226
rect 493094 28170 493150 28226
rect 493218 28170 493274 28226
rect 493342 28170 493398 28226
rect 492970 28046 493026 28102
rect 493094 28046 493150 28102
rect 493218 28046 493274 28102
rect 493342 28046 493398 28102
rect 492970 27922 493026 27978
rect 493094 27922 493150 27978
rect 493218 27922 493274 27978
rect 493342 27922 493398 27978
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 507250 526294 507306 526350
rect 507374 526294 507430 526350
rect 507498 526294 507554 526350
rect 507622 526294 507678 526350
rect 507250 526170 507306 526226
rect 507374 526170 507430 526226
rect 507498 526170 507554 526226
rect 507622 526170 507678 526226
rect 507250 526046 507306 526102
rect 507374 526046 507430 526102
rect 507498 526046 507554 526102
rect 507622 526046 507678 526102
rect 507250 525922 507306 525978
rect 507374 525922 507430 525978
rect 507498 525922 507554 525978
rect 507622 525922 507678 525978
rect 507250 508294 507306 508350
rect 507374 508294 507430 508350
rect 507498 508294 507554 508350
rect 507622 508294 507678 508350
rect 507250 508170 507306 508226
rect 507374 508170 507430 508226
rect 507498 508170 507554 508226
rect 507622 508170 507678 508226
rect 507250 508046 507306 508102
rect 507374 508046 507430 508102
rect 507498 508046 507554 508102
rect 507622 508046 507678 508102
rect 507250 507922 507306 507978
rect 507374 507922 507430 507978
rect 507498 507922 507554 507978
rect 507622 507922 507678 507978
rect 507250 490294 507306 490350
rect 507374 490294 507430 490350
rect 507498 490294 507554 490350
rect 507622 490294 507678 490350
rect 507250 490170 507306 490226
rect 507374 490170 507430 490226
rect 507498 490170 507554 490226
rect 507622 490170 507678 490226
rect 507250 490046 507306 490102
rect 507374 490046 507430 490102
rect 507498 490046 507554 490102
rect 507622 490046 507678 490102
rect 507250 489922 507306 489978
rect 507374 489922 507430 489978
rect 507498 489922 507554 489978
rect 507622 489922 507678 489978
rect 507250 472294 507306 472350
rect 507374 472294 507430 472350
rect 507498 472294 507554 472350
rect 507622 472294 507678 472350
rect 507250 472170 507306 472226
rect 507374 472170 507430 472226
rect 507498 472170 507554 472226
rect 507622 472170 507678 472226
rect 507250 472046 507306 472102
rect 507374 472046 507430 472102
rect 507498 472046 507554 472102
rect 507622 472046 507678 472102
rect 507250 471922 507306 471978
rect 507374 471922 507430 471978
rect 507498 471922 507554 471978
rect 507622 471922 507678 471978
rect 507250 454294 507306 454350
rect 507374 454294 507430 454350
rect 507498 454294 507554 454350
rect 507622 454294 507678 454350
rect 507250 454170 507306 454226
rect 507374 454170 507430 454226
rect 507498 454170 507554 454226
rect 507622 454170 507678 454226
rect 507250 454046 507306 454102
rect 507374 454046 507430 454102
rect 507498 454046 507554 454102
rect 507622 454046 507678 454102
rect 507250 453922 507306 453978
rect 507374 453922 507430 453978
rect 507498 453922 507554 453978
rect 507622 453922 507678 453978
rect 507250 436294 507306 436350
rect 507374 436294 507430 436350
rect 507498 436294 507554 436350
rect 507622 436294 507678 436350
rect 507250 436170 507306 436226
rect 507374 436170 507430 436226
rect 507498 436170 507554 436226
rect 507622 436170 507678 436226
rect 507250 436046 507306 436102
rect 507374 436046 507430 436102
rect 507498 436046 507554 436102
rect 507622 436046 507678 436102
rect 507250 435922 507306 435978
rect 507374 435922 507430 435978
rect 507498 435922 507554 435978
rect 507622 435922 507678 435978
rect 507250 418294 507306 418350
rect 507374 418294 507430 418350
rect 507498 418294 507554 418350
rect 507622 418294 507678 418350
rect 507250 418170 507306 418226
rect 507374 418170 507430 418226
rect 507498 418170 507554 418226
rect 507622 418170 507678 418226
rect 507250 418046 507306 418102
rect 507374 418046 507430 418102
rect 507498 418046 507554 418102
rect 507622 418046 507678 418102
rect 507250 417922 507306 417978
rect 507374 417922 507430 417978
rect 507498 417922 507554 417978
rect 507622 417922 507678 417978
rect 507250 400294 507306 400350
rect 507374 400294 507430 400350
rect 507498 400294 507554 400350
rect 507622 400294 507678 400350
rect 507250 400170 507306 400226
rect 507374 400170 507430 400226
rect 507498 400170 507554 400226
rect 507622 400170 507678 400226
rect 507250 400046 507306 400102
rect 507374 400046 507430 400102
rect 507498 400046 507554 400102
rect 507622 400046 507678 400102
rect 507250 399922 507306 399978
rect 507374 399922 507430 399978
rect 507498 399922 507554 399978
rect 507622 399922 507678 399978
rect 507250 382294 507306 382350
rect 507374 382294 507430 382350
rect 507498 382294 507554 382350
rect 507622 382294 507678 382350
rect 507250 382170 507306 382226
rect 507374 382170 507430 382226
rect 507498 382170 507554 382226
rect 507622 382170 507678 382226
rect 507250 382046 507306 382102
rect 507374 382046 507430 382102
rect 507498 382046 507554 382102
rect 507622 382046 507678 382102
rect 507250 381922 507306 381978
rect 507374 381922 507430 381978
rect 507498 381922 507554 381978
rect 507622 381922 507678 381978
rect 507250 364294 507306 364350
rect 507374 364294 507430 364350
rect 507498 364294 507554 364350
rect 507622 364294 507678 364350
rect 507250 364170 507306 364226
rect 507374 364170 507430 364226
rect 507498 364170 507554 364226
rect 507622 364170 507678 364226
rect 507250 364046 507306 364102
rect 507374 364046 507430 364102
rect 507498 364046 507554 364102
rect 507622 364046 507678 364102
rect 507250 363922 507306 363978
rect 507374 363922 507430 363978
rect 507498 363922 507554 363978
rect 507622 363922 507678 363978
rect 507250 346294 507306 346350
rect 507374 346294 507430 346350
rect 507498 346294 507554 346350
rect 507622 346294 507678 346350
rect 507250 346170 507306 346226
rect 507374 346170 507430 346226
rect 507498 346170 507554 346226
rect 507622 346170 507678 346226
rect 507250 346046 507306 346102
rect 507374 346046 507430 346102
rect 507498 346046 507554 346102
rect 507622 346046 507678 346102
rect 507250 345922 507306 345978
rect 507374 345922 507430 345978
rect 507498 345922 507554 345978
rect 507622 345922 507678 345978
rect 507250 328294 507306 328350
rect 507374 328294 507430 328350
rect 507498 328294 507554 328350
rect 507622 328294 507678 328350
rect 507250 328170 507306 328226
rect 507374 328170 507430 328226
rect 507498 328170 507554 328226
rect 507622 328170 507678 328226
rect 507250 328046 507306 328102
rect 507374 328046 507430 328102
rect 507498 328046 507554 328102
rect 507622 328046 507678 328102
rect 507250 327922 507306 327978
rect 507374 327922 507430 327978
rect 507498 327922 507554 327978
rect 507622 327922 507678 327978
rect 507250 310294 507306 310350
rect 507374 310294 507430 310350
rect 507498 310294 507554 310350
rect 507622 310294 507678 310350
rect 507250 310170 507306 310226
rect 507374 310170 507430 310226
rect 507498 310170 507554 310226
rect 507622 310170 507678 310226
rect 507250 310046 507306 310102
rect 507374 310046 507430 310102
rect 507498 310046 507554 310102
rect 507622 310046 507678 310102
rect 507250 309922 507306 309978
rect 507374 309922 507430 309978
rect 507498 309922 507554 309978
rect 507622 309922 507678 309978
rect 507250 292294 507306 292350
rect 507374 292294 507430 292350
rect 507498 292294 507554 292350
rect 507622 292294 507678 292350
rect 507250 292170 507306 292226
rect 507374 292170 507430 292226
rect 507498 292170 507554 292226
rect 507622 292170 507678 292226
rect 507250 292046 507306 292102
rect 507374 292046 507430 292102
rect 507498 292046 507554 292102
rect 507622 292046 507678 292102
rect 507250 291922 507306 291978
rect 507374 291922 507430 291978
rect 507498 291922 507554 291978
rect 507622 291922 507678 291978
rect 507250 274294 507306 274350
rect 507374 274294 507430 274350
rect 507498 274294 507554 274350
rect 507622 274294 507678 274350
rect 507250 274170 507306 274226
rect 507374 274170 507430 274226
rect 507498 274170 507554 274226
rect 507622 274170 507678 274226
rect 507250 274046 507306 274102
rect 507374 274046 507430 274102
rect 507498 274046 507554 274102
rect 507622 274046 507678 274102
rect 507250 273922 507306 273978
rect 507374 273922 507430 273978
rect 507498 273922 507554 273978
rect 507622 273922 507678 273978
rect 507250 256294 507306 256350
rect 507374 256294 507430 256350
rect 507498 256294 507554 256350
rect 507622 256294 507678 256350
rect 507250 256170 507306 256226
rect 507374 256170 507430 256226
rect 507498 256170 507554 256226
rect 507622 256170 507678 256226
rect 507250 256046 507306 256102
rect 507374 256046 507430 256102
rect 507498 256046 507554 256102
rect 507622 256046 507678 256102
rect 507250 255922 507306 255978
rect 507374 255922 507430 255978
rect 507498 255922 507554 255978
rect 507622 255922 507678 255978
rect 507250 238294 507306 238350
rect 507374 238294 507430 238350
rect 507498 238294 507554 238350
rect 507622 238294 507678 238350
rect 507250 238170 507306 238226
rect 507374 238170 507430 238226
rect 507498 238170 507554 238226
rect 507622 238170 507678 238226
rect 507250 238046 507306 238102
rect 507374 238046 507430 238102
rect 507498 238046 507554 238102
rect 507622 238046 507678 238102
rect 507250 237922 507306 237978
rect 507374 237922 507430 237978
rect 507498 237922 507554 237978
rect 507622 237922 507678 237978
rect 507250 220294 507306 220350
rect 507374 220294 507430 220350
rect 507498 220294 507554 220350
rect 507622 220294 507678 220350
rect 507250 220170 507306 220226
rect 507374 220170 507430 220226
rect 507498 220170 507554 220226
rect 507622 220170 507678 220226
rect 507250 220046 507306 220102
rect 507374 220046 507430 220102
rect 507498 220046 507554 220102
rect 507622 220046 507678 220102
rect 507250 219922 507306 219978
rect 507374 219922 507430 219978
rect 507498 219922 507554 219978
rect 507622 219922 507678 219978
rect 507250 202294 507306 202350
rect 507374 202294 507430 202350
rect 507498 202294 507554 202350
rect 507622 202294 507678 202350
rect 507250 202170 507306 202226
rect 507374 202170 507430 202226
rect 507498 202170 507554 202226
rect 507622 202170 507678 202226
rect 507250 202046 507306 202102
rect 507374 202046 507430 202102
rect 507498 202046 507554 202102
rect 507622 202046 507678 202102
rect 507250 201922 507306 201978
rect 507374 201922 507430 201978
rect 507498 201922 507554 201978
rect 507622 201922 507678 201978
rect 507250 184294 507306 184350
rect 507374 184294 507430 184350
rect 507498 184294 507554 184350
rect 507622 184294 507678 184350
rect 507250 184170 507306 184226
rect 507374 184170 507430 184226
rect 507498 184170 507554 184226
rect 507622 184170 507678 184226
rect 507250 184046 507306 184102
rect 507374 184046 507430 184102
rect 507498 184046 507554 184102
rect 507622 184046 507678 184102
rect 507250 183922 507306 183978
rect 507374 183922 507430 183978
rect 507498 183922 507554 183978
rect 507622 183922 507678 183978
rect 507250 166294 507306 166350
rect 507374 166294 507430 166350
rect 507498 166294 507554 166350
rect 507622 166294 507678 166350
rect 507250 166170 507306 166226
rect 507374 166170 507430 166226
rect 507498 166170 507554 166226
rect 507622 166170 507678 166226
rect 507250 166046 507306 166102
rect 507374 166046 507430 166102
rect 507498 166046 507554 166102
rect 507622 166046 507678 166102
rect 507250 165922 507306 165978
rect 507374 165922 507430 165978
rect 507498 165922 507554 165978
rect 507622 165922 507678 165978
rect 507250 148294 507306 148350
rect 507374 148294 507430 148350
rect 507498 148294 507554 148350
rect 507622 148294 507678 148350
rect 507250 148170 507306 148226
rect 507374 148170 507430 148226
rect 507498 148170 507554 148226
rect 507622 148170 507678 148226
rect 507250 148046 507306 148102
rect 507374 148046 507430 148102
rect 507498 148046 507554 148102
rect 507622 148046 507678 148102
rect 507250 147922 507306 147978
rect 507374 147922 507430 147978
rect 507498 147922 507554 147978
rect 507622 147922 507678 147978
rect 507250 130294 507306 130350
rect 507374 130294 507430 130350
rect 507498 130294 507554 130350
rect 507622 130294 507678 130350
rect 507250 130170 507306 130226
rect 507374 130170 507430 130226
rect 507498 130170 507554 130226
rect 507622 130170 507678 130226
rect 507250 130046 507306 130102
rect 507374 130046 507430 130102
rect 507498 130046 507554 130102
rect 507622 130046 507678 130102
rect 507250 129922 507306 129978
rect 507374 129922 507430 129978
rect 507498 129922 507554 129978
rect 507622 129922 507678 129978
rect 507250 112294 507306 112350
rect 507374 112294 507430 112350
rect 507498 112294 507554 112350
rect 507622 112294 507678 112350
rect 507250 112170 507306 112226
rect 507374 112170 507430 112226
rect 507498 112170 507554 112226
rect 507622 112170 507678 112226
rect 507250 112046 507306 112102
rect 507374 112046 507430 112102
rect 507498 112046 507554 112102
rect 507622 112046 507678 112102
rect 507250 111922 507306 111978
rect 507374 111922 507430 111978
rect 507498 111922 507554 111978
rect 507622 111922 507678 111978
rect 507250 94294 507306 94350
rect 507374 94294 507430 94350
rect 507498 94294 507554 94350
rect 507622 94294 507678 94350
rect 507250 94170 507306 94226
rect 507374 94170 507430 94226
rect 507498 94170 507554 94226
rect 507622 94170 507678 94226
rect 507250 94046 507306 94102
rect 507374 94046 507430 94102
rect 507498 94046 507554 94102
rect 507622 94046 507678 94102
rect 507250 93922 507306 93978
rect 507374 93922 507430 93978
rect 507498 93922 507554 93978
rect 507622 93922 507678 93978
rect 507250 76294 507306 76350
rect 507374 76294 507430 76350
rect 507498 76294 507554 76350
rect 507622 76294 507678 76350
rect 507250 76170 507306 76226
rect 507374 76170 507430 76226
rect 507498 76170 507554 76226
rect 507622 76170 507678 76226
rect 507250 76046 507306 76102
rect 507374 76046 507430 76102
rect 507498 76046 507554 76102
rect 507622 76046 507678 76102
rect 507250 75922 507306 75978
rect 507374 75922 507430 75978
rect 507498 75922 507554 75978
rect 507622 75922 507678 75978
rect 507250 58294 507306 58350
rect 507374 58294 507430 58350
rect 507498 58294 507554 58350
rect 507622 58294 507678 58350
rect 507250 58170 507306 58226
rect 507374 58170 507430 58226
rect 507498 58170 507554 58226
rect 507622 58170 507678 58226
rect 507250 58046 507306 58102
rect 507374 58046 507430 58102
rect 507498 58046 507554 58102
rect 507622 58046 507678 58102
rect 507250 57922 507306 57978
rect 507374 57922 507430 57978
rect 507498 57922 507554 57978
rect 507622 57922 507678 57978
rect 507250 40294 507306 40350
rect 507374 40294 507430 40350
rect 507498 40294 507554 40350
rect 507622 40294 507678 40350
rect 507250 40170 507306 40226
rect 507374 40170 507430 40226
rect 507498 40170 507554 40226
rect 507622 40170 507678 40226
rect 507250 40046 507306 40102
rect 507374 40046 507430 40102
rect 507498 40046 507554 40102
rect 507622 40046 507678 40102
rect 507250 39922 507306 39978
rect 507374 39922 507430 39978
rect 507498 39922 507554 39978
rect 507622 39922 507678 39978
rect 507250 22294 507306 22350
rect 507374 22294 507430 22350
rect 507498 22294 507554 22350
rect 507622 22294 507678 22350
rect 507250 22170 507306 22226
rect 507374 22170 507430 22226
rect 507498 22170 507554 22226
rect 507622 22170 507678 22226
rect 507250 22046 507306 22102
rect 507374 22046 507430 22102
rect 507498 22046 507554 22102
rect 507622 22046 507678 22102
rect 507250 21922 507306 21978
rect 507374 21922 507430 21978
rect 507498 21922 507554 21978
rect 507622 21922 507678 21978
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 510970 514294 511026 514350
rect 511094 514294 511150 514350
rect 511218 514294 511274 514350
rect 511342 514294 511398 514350
rect 510970 514170 511026 514226
rect 511094 514170 511150 514226
rect 511218 514170 511274 514226
rect 511342 514170 511398 514226
rect 510970 514046 511026 514102
rect 511094 514046 511150 514102
rect 511218 514046 511274 514102
rect 511342 514046 511398 514102
rect 510970 513922 511026 513978
rect 511094 513922 511150 513978
rect 511218 513922 511274 513978
rect 511342 513922 511398 513978
rect 510970 496294 511026 496350
rect 511094 496294 511150 496350
rect 511218 496294 511274 496350
rect 511342 496294 511398 496350
rect 510970 496170 511026 496226
rect 511094 496170 511150 496226
rect 511218 496170 511274 496226
rect 511342 496170 511398 496226
rect 510970 496046 511026 496102
rect 511094 496046 511150 496102
rect 511218 496046 511274 496102
rect 511342 496046 511398 496102
rect 510970 495922 511026 495978
rect 511094 495922 511150 495978
rect 511218 495922 511274 495978
rect 511342 495922 511398 495978
rect 510970 478294 511026 478350
rect 511094 478294 511150 478350
rect 511218 478294 511274 478350
rect 511342 478294 511398 478350
rect 510970 478170 511026 478226
rect 511094 478170 511150 478226
rect 511218 478170 511274 478226
rect 511342 478170 511398 478226
rect 510970 478046 511026 478102
rect 511094 478046 511150 478102
rect 511218 478046 511274 478102
rect 511342 478046 511398 478102
rect 510970 477922 511026 477978
rect 511094 477922 511150 477978
rect 511218 477922 511274 477978
rect 511342 477922 511398 477978
rect 510970 460294 511026 460350
rect 511094 460294 511150 460350
rect 511218 460294 511274 460350
rect 511342 460294 511398 460350
rect 510970 460170 511026 460226
rect 511094 460170 511150 460226
rect 511218 460170 511274 460226
rect 511342 460170 511398 460226
rect 510970 460046 511026 460102
rect 511094 460046 511150 460102
rect 511218 460046 511274 460102
rect 511342 460046 511398 460102
rect 510970 459922 511026 459978
rect 511094 459922 511150 459978
rect 511218 459922 511274 459978
rect 511342 459922 511398 459978
rect 510970 442294 511026 442350
rect 511094 442294 511150 442350
rect 511218 442294 511274 442350
rect 511342 442294 511398 442350
rect 510970 442170 511026 442226
rect 511094 442170 511150 442226
rect 511218 442170 511274 442226
rect 511342 442170 511398 442226
rect 510970 442046 511026 442102
rect 511094 442046 511150 442102
rect 511218 442046 511274 442102
rect 511342 442046 511398 442102
rect 510970 441922 511026 441978
rect 511094 441922 511150 441978
rect 511218 441922 511274 441978
rect 511342 441922 511398 441978
rect 510970 424294 511026 424350
rect 511094 424294 511150 424350
rect 511218 424294 511274 424350
rect 511342 424294 511398 424350
rect 510970 424170 511026 424226
rect 511094 424170 511150 424226
rect 511218 424170 511274 424226
rect 511342 424170 511398 424226
rect 510970 424046 511026 424102
rect 511094 424046 511150 424102
rect 511218 424046 511274 424102
rect 511342 424046 511398 424102
rect 510970 423922 511026 423978
rect 511094 423922 511150 423978
rect 511218 423922 511274 423978
rect 511342 423922 511398 423978
rect 510970 406294 511026 406350
rect 511094 406294 511150 406350
rect 511218 406294 511274 406350
rect 511342 406294 511398 406350
rect 510970 406170 511026 406226
rect 511094 406170 511150 406226
rect 511218 406170 511274 406226
rect 511342 406170 511398 406226
rect 510970 406046 511026 406102
rect 511094 406046 511150 406102
rect 511218 406046 511274 406102
rect 511342 406046 511398 406102
rect 510970 405922 511026 405978
rect 511094 405922 511150 405978
rect 511218 405922 511274 405978
rect 511342 405922 511398 405978
rect 510970 388294 511026 388350
rect 511094 388294 511150 388350
rect 511218 388294 511274 388350
rect 511342 388294 511398 388350
rect 510970 388170 511026 388226
rect 511094 388170 511150 388226
rect 511218 388170 511274 388226
rect 511342 388170 511398 388226
rect 510970 388046 511026 388102
rect 511094 388046 511150 388102
rect 511218 388046 511274 388102
rect 511342 388046 511398 388102
rect 510970 387922 511026 387978
rect 511094 387922 511150 387978
rect 511218 387922 511274 387978
rect 511342 387922 511398 387978
rect 510970 370294 511026 370350
rect 511094 370294 511150 370350
rect 511218 370294 511274 370350
rect 511342 370294 511398 370350
rect 510970 370170 511026 370226
rect 511094 370170 511150 370226
rect 511218 370170 511274 370226
rect 511342 370170 511398 370226
rect 510970 370046 511026 370102
rect 511094 370046 511150 370102
rect 511218 370046 511274 370102
rect 511342 370046 511398 370102
rect 510970 369922 511026 369978
rect 511094 369922 511150 369978
rect 511218 369922 511274 369978
rect 511342 369922 511398 369978
rect 510970 352294 511026 352350
rect 511094 352294 511150 352350
rect 511218 352294 511274 352350
rect 511342 352294 511398 352350
rect 510970 352170 511026 352226
rect 511094 352170 511150 352226
rect 511218 352170 511274 352226
rect 511342 352170 511398 352226
rect 510970 352046 511026 352102
rect 511094 352046 511150 352102
rect 511218 352046 511274 352102
rect 511342 352046 511398 352102
rect 510970 351922 511026 351978
rect 511094 351922 511150 351978
rect 511218 351922 511274 351978
rect 511342 351922 511398 351978
rect 510970 334294 511026 334350
rect 511094 334294 511150 334350
rect 511218 334294 511274 334350
rect 511342 334294 511398 334350
rect 510970 334170 511026 334226
rect 511094 334170 511150 334226
rect 511218 334170 511274 334226
rect 511342 334170 511398 334226
rect 510970 334046 511026 334102
rect 511094 334046 511150 334102
rect 511218 334046 511274 334102
rect 511342 334046 511398 334102
rect 510970 333922 511026 333978
rect 511094 333922 511150 333978
rect 511218 333922 511274 333978
rect 511342 333922 511398 333978
rect 510970 316294 511026 316350
rect 511094 316294 511150 316350
rect 511218 316294 511274 316350
rect 511342 316294 511398 316350
rect 510970 316170 511026 316226
rect 511094 316170 511150 316226
rect 511218 316170 511274 316226
rect 511342 316170 511398 316226
rect 510970 316046 511026 316102
rect 511094 316046 511150 316102
rect 511218 316046 511274 316102
rect 511342 316046 511398 316102
rect 510970 315922 511026 315978
rect 511094 315922 511150 315978
rect 511218 315922 511274 315978
rect 511342 315922 511398 315978
rect 510970 298294 511026 298350
rect 511094 298294 511150 298350
rect 511218 298294 511274 298350
rect 511342 298294 511398 298350
rect 510970 298170 511026 298226
rect 511094 298170 511150 298226
rect 511218 298170 511274 298226
rect 511342 298170 511398 298226
rect 510970 298046 511026 298102
rect 511094 298046 511150 298102
rect 511218 298046 511274 298102
rect 511342 298046 511398 298102
rect 510970 297922 511026 297978
rect 511094 297922 511150 297978
rect 511218 297922 511274 297978
rect 511342 297922 511398 297978
rect 510970 280294 511026 280350
rect 511094 280294 511150 280350
rect 511218 280294 511274 280350
rect 511342 280294 511398 280350
rect 510970 280170 511026 280226
rect 511094 280170 511150 280226
rect 511218 280170 511274 280226
rect 511342 280170 511398 280226
rect 510970 280046 511026 280102
rect 511094 280046 511150 280102
rect 511218 280046 511274 280102
rect 511342 280046 511398 280102
rect 510970 279922 511026 279978
rect 511094 279922 511150 279978
rect 511218 279922 511274 279978
rect 511342 279922 511398 279978
rect 510970 262294 511026 262350
rect 511094 262294 511150 262350
rect 511218 262294 511274 262350
rect 511342 262294 511398 262350
rect 510970 262170 511026 262226
rect 511094 262170 511150 262226
rect 511218 262170 511274 262226
rect 511342 262170 511398 262226
rect 510970 262046 511026 262102
rect 511094 262046 511150 262102
rect 511218 262046 511274 262102
rect 511342 262046 511398 262102
rect 510970 261922 511026 261978
rect 511094 261922 511150 261978
rect 511218 261922 511274 261978
rect 511342 261922 511398 261978
rect 510970 244294 511026 244350
rect 511094 244294 511150 244350
rect 511218 244294 511274 244350
rect 511342 244294 511398 244350
rect 510970 244170 511026 244226
rect 511094 244170 511150 244226
rect 511218 244170 511274 244226
rect 511342 244170 511398 244226
rect 510970 244046 511026 244102
rect 511094 244046 511150 244102
rect 511218 244046 511274 244102
rect 511342 244046 511398 244102
rect 510970 243922 511026 243978
rect 511094 243922 511150 243978
rect 511218 243922 511274 243978
rect 511342 243922 511398 243978
rect 510970 226294 511026 226350
rect 511094 226294 511150 226350
rect 511218 226294 511274 226350
rect 511342 226294 511398 226350
rect 510970 226170 511026 226226
rect 511094 226170 511150 226226
rect 511218 226170 511274 226226
rect 511342 226170 511398 226226
rect 510970 226046 511026 226102
rect 511094 226046 511150 226102
rect 511218 226046 511274 226102
rect 511342 226046 511398 226102
rect 510970 225922 511026 225978
rect 511094 225922 511150 225978
rect 511218 225922 511274 225978
rect 511342 225922 511398 225978
rect 510970 208294 511026 208350
rect 511094 208294 511150 208350
rect 511218 208294 511274 208350
rect 511342 208294 511398 208350
rect 510970 208170 511026 208226
rect 511094 208170 511150 208226
rect 511218 208170 511274 208226
rect 511342 208170 511398 208226
rect 510970 208046 511026 208102
rect 511094 208046 511150 208102
rect 511218 208046 511274 208102
rect 511342 208046 511398 208102
rect 510970 207922 511026 207978
rect 511094 207922 511150 207978
rect 511218 207922 511274 207978
rect 511342 207922 511398 207978
rect 510970 190294 511026 190350
rect 511094 190294 511150 190350
rect 511218 190294 511274 190350
rect 511342 190294 511398 190350
rect 510970 190170 511026 190226
rect 511094 190170 511150 190226
rect 511218 190170 511274 190226
rect 511342 190170 511398 190226
rect 510970 190046 511026 190102
rect 511094 190046 511150 190102
rect 511218 190046 511274 190102
rect 511342 190046 511398 190102
rect 510970 189922 511026 189978
rect 511094 189922 511150 189978
rect 511218 189922 511274 189978
rect 511342 189922 511398 189978
rect 510970 172294 511026 172350
rect 511094 172294 511150 172350
rect 511218 172294 511274 172350
rect 511342 172294 511398 172350
rect 510970 172170 511026 172226
rect 511094 172170 511150 172226
rect 511218 172170 511274 172226
rect 511342 172170 511398 172226
rect 510970 172046 511026 172102
rect 511094 172046 511150 172102
rect 511218 172046 511274 172102
rect 511342 172046 511398 172102
rect 510970 171922 511026 171978
rect 511094 171922 511150 171978
rect 511218 171922 511274 171978
rect 511342 171922 511398 171978
rect 510970 154294 511026 154350
rect 511094 154294 511150 154350
rect 511218 154294 511274 154350
rect 511342 154294 511398 154350
rect 510970 154170 511026 154226
rect 511094 154170 511150 154226
rect 511218 154170 511274 154226
rect 511342 154170 511398 154226
rect 510970 154046 511026 154102
rect 511094 154046 511150 154102
rect 511218 154046 511274 154102
rect 511342 154046 511398 154102
rect 510970 153922 511026 153978
rect 511094 153922 511150 153978
rect 511218 153922 511274 153978
rect 511342 153922 511398 153978
rect 510970 136294 511026 136350
rect 511094 136294 511150 136350
rect 511218 136294 511274 136350
rect 511342 136294 511398 136350
rect 510970 136170 511026 136226
rect 511094 136170 511150 136226
rect 511218 136170 511274 136226
rect 511342 136170 511398 136226
rect 510970 136046 511026 136102
rect 511094 136046 511150 136102
rect 511218 136046 511274 136102
rect 511342 136046 511398 136102
rect 510970 135922 511026 135978
rect 511094 135922 511150 135978
rect 511218 135922 511274 135978
rect 511342 135922 511398 135978
rect 510970 118294 511026 118350
rect 511094 118294 511150 118350
rect 511218 118294 511274 118350
rect 511342 118294 511398 118350
rect 510970 118170 511026 118226
rect 511094 118170 511150 118226
rect 511218 118170 511274 118226
rect 511342 118170 511398 118226
rect 510970 118046 511026 118102
rect 511094 118046 511150 118102
rect 511218 118046 511274 118102
rect 511342 118046 511398 118102
rect 510970 117922 511026 117978
rect 511094 117922 511150 117978
rect 511218 117922 511274 117978
rect 511342 117922 511398 117978
rect 510970 100294 511026 100350
rect 511094 100294 511150 100350
rect 511218 100294 511274 100350
rect 511342 100294 511398 100350
rect 510970 100170 511026 100226
rect 511094 100170 511150 100226
rect 511218 100170 511274 100226
rect 511342 100170 511398 100226
rect 510970 100046 511026 100102
rect 511094 100046 511150 100102
rect 511218 100046 511274 100102
rect 511342 100046 511398 100102
rect 510970 99922 511026 99978
rect 511094 99922 511150 99978
rect 511218 99922 511274 99978
rect 511342 99922 511398 99978
rect 510970 82294 511026 82350
rect 511094 82294 511150 82350
rect 511218 82294 511274 82350
rect 511342 82294 511398 82350
rect 510970 82170 511026 82226
rect 511094 82170 511150 82226
rect 511218 82170 511274 82226
rect 511342 82170 511398 82226
rect 510970 82046 511026 82102
rect 511094 82046 511150 82102
rect 511218 82046 511274 82102
rect 511342 82046 511398 82102
rect 510970 81922 511026 81978
rect 511094 81922 511150 81978
rect 511218 81922 511274 81978
rect 511342 81922 511398 81978
rect 510970 64294 511026 64350
rect 511094 64294 511150 64350
rect 511218 64294 511274 64350
rect 511342 64294 511398 64350
rect 510970 64170 511026 64226
rect 511094 64170 511150 64226
rect 511218 64170 511274 64226
rect 511342 64170 511398 64226
rect 510970 64046 511026 64102
rect 511094 64046 511150 64102
rect 511218 64046 511274 64102
rect 511342 64046 511398 64102
rect 510970 63922 511026 63978
rect 511094 63922 511150 63978
rect 511218 63922 511274 63978
rect 511342 63922 511398 63978
rect 510970 46294 511026 46350
rect 511094 46294 511150 46350
rect 511218 46294 511274 46350
rect 511342 46294 511398 46350
rect 510970 46170 511026 46226
rect 511094 46170 511150 46226
rect 511218 46170 511274 46226
rect 511342 46170 511398 46226
rect 510970 46046 511026 46102
rect 511094 46046 511150 46102
rect 511218 46046 511274 46102
rect 511342 46046 511398 46102
rect 510970 45922 511026 45978
rect 511094 45922 511150 45978
rect 511218 45922 511274 45978
rect 511342 45922 511398 45978
rect 510970 28294 511026 28350
rect 511094 28294 511150 28350
rect 511218 28294 511274 28350
rect 511342 28294 511398 28350
rect 510970 28170 511026 28226
rect 511094 28170 511150 28226
rect 511218 28170 511274 28226
rect 511342 28170 511398 28226
rect 510970 28046 511026 28102
rect 511094 28046 511150 28102
rect 511218 28046 511274 28102
rect 511342 28046 511398 28102
rect 510970 27922 511026 27978
rect 511094 27922 511150 27978
rect 511218 27922 511274 27978
rect 511342 27922 511398 27978
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 525250 597156 525306 597212
rect 525374 597156 525430 597212
rect 525498 597156 525554 597212
rect 525622 597156 525678 597212
rect 525250 597032 525306 597088
rect 525374 597032 525430 597088
rect 525498 597032 525554 597088
rect 525622 597032 525678 597088
rect 525250 596908 525306 596964
rect 525374 596908 525430 596964
rect 525498 596908 525554 596964
rect 525622 596908 525678 596964
rect 525250 596784 525306 596840
rect 525374 596784 525430 596840
rect 525498 596784 525554 596840
rect 525622 596784 525678 596840
rect 525250 580294 525306 580350
rect 525374 580294 525430 580350
rect 525498 580294 525554 580350
rect 525622 580294 525678 580350
rect 525250 580170 525306 580226
rect 525374 580170 525430 580226
rect 525498 580170 525554 580226
rect 525622 580170 525678 580226
rect 525250 580046 525306 580102
rect 525374 580046 525430 580102
rect 525498 580046 525554 580102
rect 525622 580046 525678 580102
rect 525250 579922 525306 579978
rect 525374 579922 525430 579978
rect 525498 579922 525554 579978
rect 525622 579922 525678 579978
rect 525250 562294 525306 562350
rect 525374 562294 525430 562350
rect 525498 562294 525554 562350
rect 525622 562294 525678 562350
rect 525250 562170 525306 562226
rect 525374 562170 525430 562226
rect 525498 562170 525554 562226
rect 525622 562170 525678 562226
rect 525250 562046 525306 562102
rect 525374 562046 525430 562102
rect 525498 562046 525554 562102
rect 525622 562046 525678 562102
rect 525250 561922 525306 561978
rect 525374 561922 525430 561978
rect 525498 561922 525554 561978
rect 525622 561922 525678 561978
rect 525250 544294 525306 544350
rect 525374 544294 525430 544350
rect 525498 544294 525554 544350
rect 525622 544294 525678 544350
rect 525250 544170 525306 544226
rect 525374 544170 525430 544226
rect 525498 544170 525554 544226
rect 525622 544170 525678 544226
rect 525250 544046 525306 544102
rect 525374 544046 525430 544102
rect 525498 544046 525554 544102
rect 525622 544046 525678 544102
rect 525250 543922 525306 543978
rect 525374 543922 525430 543978
rect 525498 543922 525554 543978
rect 525622 543922 525678 543978
rect 525250 526294 525306 526350
rect 525374 526294 525430 526350
rect 525498 526294 525554 526350
rect 525622 526294 525678 526350
rect 525250 526170 525306 526226
rect 525374 526170 525430 526226
rect 525498 526170 525554 526226
rect 525622 526170 525678 526226
rect 525250 526046 525306 526102
rect 525374 526046 525430 526102
rect 525498 526046 525554 526102
rect 525622 526046 525678 526102
rect 525250 525922 525306 525978
rect 525374 525922 525430 525978
rect 525498 525922 525554 525978
rect 525622 525922 525678 525978
rect 525250 508294 525306 508350
rect 525374 508294 525430 508350
rect 525498 508294 525554 508350
rect 525622 508294 525678 508350
rect 525250 508170 525306 508226
rect 525374 508170 525430 508226
rect 525498 508170 525554 508226
rect 525622 508170 525678 508226
rect 525250 508046 525306 508102
rect 525374 508046 525430 508102
rect 525498 508046 525554 508102
rect 525622 508046 525678 508102
rect 525250 507922 525306 507978
rect 525374 507922 525430 507978
rect 525498 507922 525554 507978
rect 525622 507922 525678 507978
rect 525250 490294 525306 490350
rect 525374 490294 525430 490350
rect 525498 490294 525554 490350
rect 525622 490294 525678 490350
rect 525250 490170 525306 490226
rect 525374 490170 525430 490226
rect 525498 490170 525554 490226
rect 525622 490170 525678 490226
rect 525250 490046 525306 490102
rect 525374 490046 525430 490102
rect 525498 490046 525554 490102
rect 525622 490046 525678 490102
rect 525250 489922 525306 489978
rect 525374 489922 525430 489978
rect 525498 489922 525554 489978
rect 525622 489922 525678 489978
rect 525250 472294 525306 472350
rect 525374 472294 525430 472350
rect 525498 472294 525554 472350
rect 525622 472294 525678 472350
rect 525250 472170 525306 472226
rect 525374 472170 525430 472226
rect 525498 472170 525554 472226
rect 525622 472170 525678 472226
rect 525250 472046 525306 472102
rect 525374 472046 525430 472102
rect 525498 472046 525554 472102
rect 525622 472046 525678 472102
rect 525250 471922 525306 471978
rect 525374 471922 525430 471978
rect 525498 471922 525554 471978
rect 525622 471922 525678 471978
rect 525250 454294 525306 454350
rect 525374 454294 525430 454350
rect 525498 454294 525554 454350
rect 525622 454294 525678 454350
rect 525250 454170 525306 454226
rect 525374 454170 525430 454226
rect 525498 454170 525554 454226
rect 525622 454170 525678 454226
rect 525250 454046 525306 454102
rect 525374 454046 525430 454102
rect 525498 454046 525554 454102
rect 525622 454046 525678 454102
rect 525250 453922 525306 453978
rect 525374 453922 525430 453978
rect 525498 453922 525554 453978
rect 525622 453922 525678 453978
rect 525250 436294 525306 436350
rect 525374 436294 525430 436350
rect 525498 436294 525554 436350
rect 525622 436294 525678 436350
rect 525250 436170 525306 436226
rect 525374 436170 525430 436226
rect 525498 436170 525554 436226
rect 525622 436170 525678 436226
rect 525250 436046 525306 436102
rect 525374 436046 525430 436102
rect 525498 436046 525554 436102
rect 525622 436046 525678 436102
rect 525250 435922 525306 435978
rect 525374 435922 525430 435978
rect 525498 435922 525554 435978
rect 525622 435922 525678 435978
rect 525250 418294 525306 418350
rect 525374 418294 525430 418350
rect 525498 418294 525554 418350
rect 525622 418294 525678 418350
rect 525250 418170 525306 418226
rect 525374 418170 525430 418226
rect 525498 418170 525554 418226
rect 525622 418170 525678 418226
rect 525250 418046 525306 418102
rect 525374 418046 525430 418102
rect 525498 418046 525554 418102
rect 525622 418046 525678 418102
rect 525250 417922 525306 417978
rect 525374 417922 525430 417978
rect 525498 417922 525554 417978
rect 525622 417922 525678 417978
rect 525250 400294 525306 400350
rect 525374 400294 525430 400350
rect 525498 400294 525554 400350
rect 525622 400294 525678 400350
rect 525250 400170 525306 400226
rect 525374 400170 525430 400226
rect 525498 400170 525554 400226
rect 525622 400170 525678 400226
rect 525250 400046 525306 400102
rect 525374 400046 525430 400102
rect 525498 400046 525554 400102
rect 525622 400046 525678 400102
rect 525250 399922 525306 399978
rect 525374 399922 525430 399978
rect 525498 399922 525554 399978
rect 525622 399922 525678 399978
rect 525250 382294 525306 382350
rect 525374 382294 525430 382350
rect 525498 382294 525554 382350
rect 525622 382294 525678 382350
rect 525250 382170 525306 382226
rect 525374 382170 525430 382226
rect 525498 382170 525554 382226
rect 525622 382170 525678 382226
rect 525250 382046 525306 382102
rect 525374 382046 525430 382102
rect 525498 382046 525554 382102
rect 525622 382046 525678 382102
rect 525250 381922 525306 381978
rect 525374 381922 525430 381978
rect 525498 381922 525554 381978
rect 525622 381922 525678 381978
rect 525250 364294 525306 364350
rect 525374 364294 525430 364350
rect 525498 364294 525554 364350
rect 525622 364294 525678 364350
rect 525250 364170 525306 364226
rect 525374 364170 525430 364226
rect 525498 364170 525554 364226
rect 525622 364170 525678 364226
rect 525250 364046 525306 364102
rect 525374 364046 525430 364102
rect 525498 364046 525554 364102
rect 525622 364046 525678 364102
rect 525250 363922 525306 363978
rect 525374 363922 525430 363978
rect 525498 363922 525554 363978
rect 525622 363922 525678 363978
rect 525250 346294 525306 346350
rect 525374 346294 525430 346350
rect 525498 346294 525554 346350
rect 525622 346294 525678 346350
rect 525250 346170 525306 346226
rect 525374 346170 525430 346226
rect 525498 346170 525554 346226
rect 525622 346170 525678 346226
rect 525250 346046 525306 346102
rect 525374 346046 525430 346102
rect 525498 346046 525554 346102
rect 525622 346046 525678 346102
rect 525250 345922 525306 345978
rect 525374 345922 525430 345978
rect 525498 345922 525554 345978
rect 525622 345922 525678 345978
rect 525250 328294 525306 328350
rect 525374 328294 525430 328350
rect 525498 328294 525554 328350
rect 525622 328294 525678 328350
rect 525250 328170 525306 328226
rect 525374 328170 525430 328226
rect 525498 328170 525554 328226
rect 525622 328170 525678 328226
rect 525250 328046 525306 328102
rect 525374 328046 525430 328102
rect 525498 328046 525554 328102
rect 525622 328046 525678 328102
rect 525250 327922 525306 327978
rect 525374 327922 525430 327978
rect 525498 327922 525554 327978
rect 525622 327922 525678 327978
rect 525250 310294 525306 310350
rect 525374 310294 525430 310350
rect 525498 310294 525554 310350
rect 525622 310294 525678 310350
rect 525250 310170 525306 310226
rect 525374 310170 525430 310226
rect 525498 310170 525554 310226
rect 525622 310170 525678 310226
rect 525250 310046 525306 310102
rect 525374 310046 525430 310102
rect 525498 310046 525554 310102
rect 525622 310046 525678 310102
rect 525250 309922 525306 309978
rect 525374 309922 525430 309978
rect 525498 309922 525554 309978
rect 525622 309922 525678 309978
rect 525250 292294 525306 292350
rect 525374 292294 525430 292350
rect 525498 292294 525554 292350
rect 525622 292294 525678 292350
rect 525250 292170 525306 292226
rect 525374 292170 525430 292226
rect 525498 292170 525554 292226
rect 525622 292170 525678 292226
rect 525250 292046 525306 292102
rect 525374 292046 525430 292102
rect 525498 292046 525554 292102
rect 525622 292046 525678 292102
rect 525250 291922 525306 291978
rect 525374 291922 525430 291978
rect 525498 291922 525554 291978
rect 525622 291922 525678 291978
rect 525250 274294 525306 274350
rect 525374 274294 525430 274350
rect 525498 274294 525554 274350
rect 525622 274294 525678 274350
rect 525250 274170 525306 274226
rect 525374 274170 525430 274226
rect 525498 274170 525554 274226
rect 525622 274170 525678 274226
rect 525250 274046 525306 274102
rect 525374 274046 525430 274102
rect 525498 274046 525554 274102
rect 525622 274046 525678 274102
rect 525250 273922 525306 273978
rect 525374 273922 525430 273978
rect 525498 273922 525554 273978
rect 525622 273922 525678 273978
rect 525250 256294 525306 256350
rect 525374 256294 525430 256350
rect 525498 256294 525554 256350
rect 525622 256294 525678 256350
rect 525250 256170 525306 256226
rect 525374 256170 525430 256226
rect 525498 256170 525554 256226
rect 525622 256170 525678 256226
rect 525250 256046 525306 256102
rect 525374 256046 525430 256102
rect 525498 256046 525554 256102
rect 525622 256046 525678 256102
rect 525250 255922 525306 255978
rect 525374 255922 525430 255978
rect 525498 255922 525554 255978
rect 525622 255922 525678 255978
rect 525250 238294 525306 238350
rect 525374 238294 525430 238350
rect 525498 238294 525554 238350
rect 525622 238294 525678 238350
rect 525250 238170 525306 238226
rect 525374 238170 525430 238226
rect 525498 238170 525554 238226
rect 525622 238170 525678 238226
rect 525250 238046 525306 238102
rect 525374 238046 525430 238102
rect 525498 238046 525554 238102
rect 525622 238046 525678 238102
rect 525250 237922 525306 237978
rect 525374 237922 525430 237978
rect 525498 237922 525554 237978
rect 525622 237922 525678 237978
rect 525250 220294 525306 220350
rect 525374 220294 525430 220350
rect 525498 220294 525554 220350
rect 525622 220294 525678 220350
rect 525250 220170 525306 220226
rect 525374 220170 525430 220226
rect 525498 220170 525554 220226
rect 525622 220170 525678 220226
rect 525250 220046 525306 220102
rect 525374 220046 525430 220102
rect 525498 220046 525554 220102
rect 525622 220046 525678 220102
rect 525250 219922 525306 219978
rect 525374 219922 525430 219978
rect 525498 219922 525554 219978
rect 525622 219922 525678 219978
rect 525250 202294 525306 202350
rect 525374 202294 525430 202350
rect 525498 202294 525554 202350
rect 525622 202294 525678 202350
rect 525250 202170 525306 202226
rect 525374 202170 525430 202226
rect 525498 202170 525554 202226
rect 525622 202170 525678 202226
rect 525250 202046 525306 202102
rect 525374 202046 525430 202102
rect 525498 202046 525554 202102
rect 525622 202046 525678 202102
rect 525250 201922 525306 201978
rect 525374 201922 525430 201978
rect 525498 201922 525554 201978
rect 525622 201922 525678 201978
rect 525250 184294 525306 184350
rect 525374 184294 525430 184350
rect 525498 184294 525554 184350
rect 525622 184294 525678 184350
rect 525250 184170 525306 184226
rect 525374 184170 525430 184226
rect 525498 184170 525554 184226
rect 525622 184170 525678 184226
rect 525250 184046 525306 184102
rect 525374 184046 525430 184102
rect 525498 184046 525554 184102
rect 525622 184046 525678 184102
rect 525250 183922 525306 183978
rect 525374 183922 525430 183978
rect 525498 183922 525554 183978
rect 525622 183922 525678 183978
rect 525250 166294 525306 166350
rect 525374 166294 525430 166350
rect 525498 166294 525554 166350
rect 525622 166294 525678 166350
rect 525250 166170 525306 166226
rect 525374 166170 525430 166226
rect 525498 166170 525554 166226
rect 525622 166170 525678 166226
rect 525250 166046 525306 166102
rect 525374 166046 525430 166102
rect 525498 166046 525554 166102
rect 525622 166046 525678 166102
rect 525250 165922 525306 165978
rect 525374 165922 525430 165978
rect 525498 165922 525554 165978
rect 525622 165922 525678 165978
rect 525250 148294 525306 148350
rect 525374 148294 525430 148350
rect 525498 148294 525554 148350
rect 525622 148294 525678 148350
rect 525250 148170 525306 148226
rect 525374 148170 525430 148226
rect 525498 148170 525554 148226
rect 525622 148170 525678 148226
rect 525250 148046 525306 148102
rect 525374 148046 525430 148102
rect 525498 148046 525554 148102
rect 525622 148046 525678 148102
rect 525250 147922 525306 147978
rect 525374 147922 525430 147978
rect 525498 147922 525554 147978
rect 525622 147922 525678 147978
rect 525250 130294 525306 130350
rect 525374 130294 525430 130350
rect 525498 130294 525554 130350
rect 525622 130294 525678 130350
rect 525250 130170 525306 130226
rect 525374 130170 525430 130226
rect 525498 130170 525554 130226
rect 525622 130170 525678 130226
rect 525250 130046 525306 130102
rect 525374 130046 525430 130102
rect 525498 130046 525554 130102
rect 525622 130046 525678 130102
rect 525250 129922 525306 129978
rect 525374 129922 525430 129978
rect 525498 129922 525554 129978
rect 525622 129922 525678 129978
rect 525250 112294 525306 112350
rect 525374 112294 525430 112350
rect 525498 112294 525554 112350
rect 525622 112294 525678 112350
rect 525250 112170 525306 112226
rect 525374 112170 525430 112226
rect 525498 112170 525554 112226
rect 525622 112170 525678 112226
rect 525250 112046 525306 112102
rect 525374 112046 525430 112102
rect 525498 112046 525554 112102
rect 525622 112046 525678 112102
rect 525250 111922 525306 111978
rect 525374 111922 525430 111978
rect 525498 111922 525554 111978
rect 525622 111922 525678 111978
rect 525250 94294 525306 94350
rect 525374 94294 525430 94350
rect 525498 94294 525554 94350
rect 525622 94294 525678 94350
rect 525250 94170 525306 94226
rect 525374 94170 525430 94226
rect 525498 94170 525554 94226
rect 525622 94170 525678 94226
rect 525250 94046 525306 94102
rect 525374 94046 525430 94102
rect 525498 94046 525554 94102
rect 525622 94046 525678 94102
rect 525250 93922 525306 93978
rect 525374 93922 525430 93978
rect 525498 93922 525554 93978
rect 525622 93922 525678 93978
rect 525250 76294 525306 76350
rect 525374 76294 525430 76350
rect 525498 76294 525554 76350
rect 525622 76294 525678 76350
rect 525250 76170 525306 76226
rect 525374 76170 525430 76226
rect 525498 76170 525554 76226
rect 525622 76170 525678 76226
rect 525250 76046 525306 76102
rect 525374 76046 525430 76102
rect 525498 76046 525554 76102
rect 525622 76046 525678 76102
rect 525250 75922 525306 75978
rect 525374 75922 525430 75978
rect 525498 75922 525554 75978
rect 525622 75922 525678 75978
rect 525250 58294 525306 58350
rect 525374 58294 525430 58350
rect 525498 58294 525554 58350
rect 525622 58294 525678 58350
rect 525250 58170 525306 58226
rect 525374 58170 525430 58226
rect 525498 58170 525554 58226
rect 525622 58170 525678 58226
rect 525250 58046 525306 58102
rect 525374 58046 525430 58102
rect 525498 58046 525554 58102
rect 525622 58046 525678 58102
rect 525250 57922 525306 57978
rect 525374 57922 525430 57978
rect 525498 57922 525554 57978
rect 525622 57922 525678 57978
rect 525250 40294 525306 40350
rect 525374 40294 525430 40350
rect 525498 40294 525554 40350
rect 525622 40294 525678 40350
rect 525250 40170 525306 40226
rect 525374 40170 525430 40226
rect 525498 40170 525554 40226
rect 525622 40170 525678 40226
rect 525250 40046 525306 40102
rect 525374 40046 525430 40102
rect 525498 40046 525554 40102
rect 525622 40046 525678 40102
rect 525250 39922 525306 39978
rect 525374 39922 525430 39978
rect 525498 39922 525554 39978
rect 525622 39922 525678 39978
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 528970 514294 529026 514350
rect 529094 514294 529150 514350
rect 529218 514294 529274 514350
rect 529342 514294 529398 514350
rect 528970 514170 529026 514226
rect 529094 514170 529150 514226
rect 529218 514170 529274 514226
rect 529342 514170 529398 514226
rect 528970 514046 529026 514102
rect 529094 514046 529150 514102
rect 529218 514046 529274 514102
rect 529342 514046 529398 514102
rect 528970 513922 529026 513978
rect 529094 513922 529150 513978
rect 529218 513922 529274 513978
rect 529342 513922 529398 513978
rect 528970 496294 529026 496350
rect 529094 496294 529150 496350
rect 529218 496294 529274 496350
rect 529342 496294 529398 496350
rect 528970 496170 529026 496226
rect 529094 496170 529150 496226
rect 529218 496170 529274 496226
rect 529342 496170 529398 496226
rect 528970 496046 529026 496102
rect 529094 496046 529150 496102
rect 529218 496046 529274 496102
rect 529342 496046 529398 496102
rect 528970 495922 529026 495978
rect 529094 495922 529150 495978
rect 529218 495922 529274 495978
rect 529342 495922 529398 495978
rect 528970 478294 529026 478350
rect 529094 478294 529150 478350
rect 529218 478294 529274 478350
rect 529342 478294 529398 478350
rect 528970 478170 529026 478226
rect 529094 478170 529150 478226
rect 529218 478170 529274 478226
rect 529342 478170 529398 478226
rect 528970 478046 529026 478102
rect 529094 478046 529150 478102
rect 529218 478046 529274 478102
rect 529342 478046 529398 478102
rect 528970 477922 529026 477978
rect 529094 477922 529150 477978
rect 529218 477922 529274 477978
rect 529342 477922 529398 477978
rect 528970 460294 529026 460350
rect 529094 460294 529150 460350
rect 529218 460294 529274 460350
rect 529342 460294 529398 460350
rect 528970 460170 529026 460226
rect 529094 460170 529150 460226
rect 529218 460170 529274 460226
rect 529342 460170 529398 460226
rect 528970 460046 529026 460102
rect 529094 460046 529150 460102
rect 529218 460046 529274 460102
rect 529342 460046 529398 460102
rect 528970 459922 529026 459978
rect 529094 459922 529150 459978
rect 529218 459922 529274 459978
rect 529342 459922 529398 459978
rect 528970 442294 529026 442350
rect 529094 442294 529150 442350
rect 529218 442294 529274 442350
rect 529342 442294 529398 442350
rect 528970 442170 529026 442226
rect 529094 442170 529150 442226
rect 529218 442170 529274 442226
rect 529342 442170 529398 442226
rect 528970 442046 529026 442102
rect 529094 442046 529150 442102
rect 529218 442046 529274 442102
rect 529342 442046 529398 442102
rect 528970 441922 529026 441978
rect 529094 441922 529150 441978
rect 529218 441922 529274 441978
rect 529342 441922 529398 441978
rect 528970 424294 529026 424350
rect 529094 424294 529150 424350
rect 529218 424294 529274 424350
rect 529342 424294 529398 424350
rect 528970 424170 529026 424226
rect 529094 424170 529150 424226
rect 529218 424170 529274 424226
rect 529342 424170 529398 424226
rect 528970 424046 529026 424102
rect 529094 424046 529150 424102
rect 529218 424046 529274 424102
rect 529342 424046 529398 424102
rect 528970 423922 529026 423978
rect 529094 423922 529150 423978
rect 529218 423922 529274 423978
rect 529342 423922 529398 423978
rect 528970 406294 529026 406350
rect 529094 406294 529150 406350
rect 529218 406294 529274 406350
rect 529342 406294 529398 406350
rect 528970 406170 529026 406226
rect 529094 406170 529150 406226
rect 529218 406170 529274 406226
rect 529342 406170 529398 406226
rect 528970 406046 529026 406102
rect 529094 406046 529150 406102
rect 529218 406046 529274 406102
rect 529342 406046 529398 406102
rect 528970 405922 529026 405978
rect 529094 405922 529150 405978
rect 529218 405922 529274 405978
rect 529342 405922 529398 405978
rect 528970 388294 529026 388350
rect 529094 388294 529150 388350
rect 529218 388294 529274 388350
rect 529342 388294 529398 388350
rect 528970 388170 529026 388226
rect 529094 388170 529150 388226
rect 529218 388170 529274 388226
rect 529342 388170 529398 388226
rect 528970 388046 529026 388102
rect 529094 388046 529150 388102
rect 529218 388046 529274 388102
rect 529342 388046 529398 388102
rect 528970 387922 529026 387978
rect 529094 387922 529150 387978
rect 529218 387922 529274 387978
rect 529342 387922 529398 387978
rect 528970 370294 529026 370350
rect 529094 370294 529150 370350
rect 529218 370294 529274 370350
rect 529342 370294 529398 370350
rect 528970 370170 529026 370226
rect 529094 370170 529150 370226
rect 529218 370170 529274 370226
rect 529342 370170 529398 370226
rect 528970 370046 529026 370102
rect 529094 370046 529150 370102
rect 529218 370046 529274 370102
rect 529342 370046 529398 370102
rect 528970 369922 529026 369978
rect 529094 369922 529150 369978
rect 529218 369922 529274 369978
rect 529342 369922 529398 369978
rect 528970 352294 529026 352350
rect 529094 352294 529150 352350
rect 529218 352294 529274 352350
rect 529342 352294 529398 352350
rect 528970 352170 529026 352226
rect 529094 352170 529150 352226
rect 529218 352170 529274 352226
rect 529342 352170 529398 352226
rect 528970 352046 529026 352102
rect 529094 352046 529150 352102
rect 529218 352046 529274 352102
rect 529342 352046 529398 352102
rect 528970 351922 529026 351978
rect 529094 351922 529150 351978
rect 529218 351922 529274 351978
rect 529342 351922 529398 351978
rect 528970 334294 529026 334350
rect 529094 334294 529150 334350
rect 529218 334294 529274 334350
rect 529342 334294 529398 334350
rect 528970 334170 529026 334226
rect 529094 334170 529150 334226
rect 529218 334170 529274 334226
rect 529342 334170 529398 334226
rect 528970 334046 529026 334102
rect 529094 334046 529150 334102
rect 529218 334046 529274 334102
rect 529342 334046 529398 334102
rect 528970 333922 529026 333978
rect 529094 333922 529150 333978
rect 529218 333922 529274 333978
rect 529342 333922 529398 333978
rect 528970 316294 529026 316350
rect 529094 316294 529150 316350
rect 529218 316294 529274 316350
rect 529342 316294 529398 316350
rect 528970 316170 529026 316226
rect 529094 316170 529150 316226
rect 529218 316170 529274 316226
rect 529342 316170 529398 316226
rect 528970 316046 529026 316102
rect 529094 316046 529150 316102
rect 529218 316046 529274 316102
rect 529342 316046 529398 316102
rect 528970 315922 529026 315978
rect 529094 315922 529150 315978
rect 529218 315922 529274 315978
rect 529342 315922 529398 315978
rect 528970 298294 529026 298350
rect 529094 298294 529150 298350
rect 529218 298294 529274 298350
rect 529342 298294 529398 298350
rect 528970 298170 529026 298226
rect 529094 298170 529150 298226
rect 529218 298170 529274 298226
rect 529342 298170 529398 298226
rect 528970 298046 529026 298102
rect 529094 298046 529150 298102
rect 529218 298046 529274 298102
rect 529342 298046 529398 298102
rect 528970 297922 529026 297978
rect 529094 297922 529150 297978
rect 529218 297922 529274 297978
rect 529342 297922 529398 297978
rect 528970 280294 529026 280350
rect 529094 280294 529150 280350
rect 529218 280294 529274 280350
rect 529342 280294 529398 280350
rect 528970 280170 529026 280226
rect 529094 280170 529150 280226
rect 529218 280170 529274 280226
rect 529342 280170 529398 280226
rect 528970 280046 529026 280102
rect 529094 280046 529150 280102
rect 529218 280046 529274 280102
rect 529342 280046 529398 280102
rect 528970 279922 529026 279978
rect 529094 279922 529150 279978
rect 529218 279922 529274 279978
rect 529342 279922 529398 279978
rect 528970 262294 529026 262350
rect 529094 262294 529150 262350
rect 529218 262294 529274 262350
rect 529342 262294 529398 262350
rect 528970 262170 529026 262226
rect 529094 262170 529150 262226
rect 529218 262170 529274 262226
rect 529342 262170 529398 262226
rect 528970 262046 529026 262102
rect 529094 262046 529150 262102
rect 529218 262046 529274 262102
rect 529342 262046 529398 262102
rect 528970 261922 529026 261978
rect 529094 261922 529150 261978
rect 529218 261922 529274 261978
rect 529342 261922 529398 261978
rect 528970 244294 529026 244350
rect 529094 244294 529150 244350
rect 529218 244294 529274 244350
rect 529342 244294 529398 244350
rect 528970 244170 529026 244226
rect 529094 244170 529150 244226
rect 529218 244170 529274 244226
rect 529342 244170 529398 244226
rect 528970 244046 529026 244102
rect 529094 244046 529150 244102
rect 529218 244046 529274 244102
rect 529342 244046 529398 244102
rect 528970 243922 529026 243978
rect 529094 243922 529150 243978
rect 529218 243922 529274 243978
rect 529342 243922 529398 243978
rect 528970 226294 529026 226350
rect 529094 226294 529150 226350
rect 529218 226294 529274 226350
rect 529342 226294 529398 226350
rect 528970 226170 529026 226226
rect 529094 226170 529150 226226
rect 529218 226170 529274 226226
rect 529342 226170 529398 226226
rect 528970 226046 529026 226102
rect 529094 226046 529150 226102
rect 529218 226046 529274 226102
rect 529342 226046 529398 226102
rect 528970 225922 529026 225978
rect 529094 225922 529150 225978
rect 529218 225922 529274 225978
rect 529342 225922 529398 225978
rect 528970 208294 529026 208350
rect 529094 208294 529150 208350
rect 529218 208294 529274 208350
rect 529342 208294 529398 208350
rect 528970 208170 529026 208226
rect 529094 208170 529150 208226
rect 529218 208170 529274 208226
rect 529342 208170 529398 208226
rect 528970 208046 529026 208102
rect 529094 208046 529150 208102
rect 529218 208046 529274 208102
rect 529342 208046 529398 208102
rect 528970 207922 529026 207978
rect 529094 207922 529150 207978
rect 529218 207922 529274 207978
rect 529342 207922 529398 207978
rect 528970 190294 529026 190350
rect 529094 190294 529150 190350
rect 529218 190294 529274 190350
rect 529342 190294 529398 190350
rect 528970 190170 529026 190226
rect 529094 190170 529150 190226
rect 529218 190170 529274 190226
rect 529342 190170 529398 190226
rect 528970 190046 529026 190102
rect 529094 190046 529150 190102
rect 529218 190046 529274 190102
rect 529342 190046 529398 190102
rect 528970 189922 529026 189978
rect 529094 189922 529150 189978
rect 529218 189922 529274 189978
rect 529342 189922 529398 189978
rect 528970 172294 529026 172350
rect 529094 172294 529150 172350
rect 529218 172294 529274 172350
rect 529342 172294 529398 172350
rect 528970 172170 529026 172226
rect 529094 172170 529150 172226
rect 529218 172170 529274 172226
rect 529342 172170 529398 172226
rect 528970 172046 529026 172102
rect 529094 172046 529150 172102
rect 529218 172046 529274 172102
rect 529342 172046 529398 172102
rect 528970 171922 529026 171978
rect 529094 171922 529150 171978
rect 529218 171922 529274 171978
rect 529342 171922 529398 171978
rect 528970 154294 529026 154350
rect 529094 154294 529150 154350
rect 529218 154294 529274 154350
rect 529342 154294 529398 154350
rect 528970 154170 529026 154226
rect 529094 154170 529150 154226
rect 529218 154170 529274 154226
rect 529342 154170 529398 154226
rect 528970 154046 529026 154102
rect 529094 154046 529150 154102
rect 529218 154046 529274 154102
rect 529342 154046 529398 154102
rect 528970 153922 529026 153978
rect 529094 153922 529150 153978
rect 529218 153922 529274 153978
rect 529342 153922 529398 153978
rect 528970 136294 529026 136350
rect 529094 136294 529150 136350
rect 529218 136294 529274 136350
rect 529342 136294 529398 136350
rect 528970 136170 529026 136226
rect 529094 136170 529150 136226
rect 529218 136170 529274 136226
rect 529342 136170 529398 136226
rect 528970 136046 529026 136102
rect 529094 136046 529150 136102
rect 529218 136046 529274 136102
rect 529342 136046 529398 136102
rect 528970 135922 529026 135978
rect 529094 135922 529150 135978
rect 529218 135922 529274 135978
rect 529342 135922 529398 135978
rect 528970 118294 529026 118350
rect 529094 118294 529150 118350
rect 529218 118294 529274 118350
rect 529342 118294 529398 118350
rect 528970 118170 529026 118226
rect 529094 118170 529150 118226
rect 529218 118170 529274 118226
rect 529342 118170 529398 118226
rect 528970 118046 529026 118102
rect 529094 118046 529150 118102
rect 529218 118046 529274 118102
rect 529342 118046 529398 118102
rect 528970 117922 529026 117978
rect 529094 117922 529150 117978
rect 529218 117922 529274 117978
rect 529342 117922 529398 117978
rect 528970 100294 529026 100350
rect 529094 100294 529150 100350
rect 529218 100294 529274 100350
rect 529342 100294 529398 100350
rect 528970 100170 529026 100226
rect 529094 100170 529150 100226
rect 529218 100170 529274 100226
rect 529342 100170 529398 100226
rect 528970 100046 529026 100102
rect 529094 100046 529150 100102
rect 529218 100046 529274 100102
rect 529342 100046 529398 100102
rect 528970 99922 529026 99978
rect 529094 99922 529150 99978
rect 529218 99922 529274 99978
rect 529342 99922 529398 99978
rect 528970 82294 529026 82350
rect 529094 82294 529150 82350
rect 529218 82294 529274 82350
rect 529342 82294 529398 82350
rect 528970 82170 529026 82226
rect 529094 82170 529150 82226
rect 529218 82170 529274 82226
rect 529342 82170 529398 82226
rect 528970 82046 529026 82102
rect 529094 82046 529150 82102
rect 529218 82046 529274 82102
rect 529342 82046 529398 82102
rect 528970 81922 529026 81978
rect 529094 81922 529150 81978
rect 529218 81922 529274 81978
rect 529342 81922 529398 81978
rect 528970 64294 529026 64350
rect 529094 64294 529150 64350
rect 529218 64294 529274 64350
rect 529342 64294 529398 64350
rect 528970 64170 529026 64226
rect 529094 64170 529150 64226
rect 529218 64170 529274 64226
rect 529342 64170 529398 64226
rect 528970 64046 529026 64102
rect 529094 64046 529150 64102
rect 529218 64046 529274 64102
rect 529342 64046 529398 64102
rect 528970 63922 529026 63978
rect 529094 63922 529150 63978
rect 529218 63922 529274 63978
rect 529342 63922 529398 63978
rect 528970 46294 529026 46350
rect 529094 46294 529150 46350
rect 529218 46294 529274 46350
rect 529342 46294 529398 46350
rect 528970 46170 529026 46226
rect 529094 46170 529150 46226
rect 529218 46170 529274 46226
rect 529342 46170 529398 46226
rect 528970 46046 529026 46102
rect 529094 46046 529150 46102
rect 529218 46046 529274 46102
rect 529342 46046 529398 46102
rect 528970 45922 529026 45978
rect 529094 45922 529150 45978
rect 529218 45922 529274 45978
rect 529342 45922 529398 45978
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 543250 526294 543306 526350
rect 543374 526294 543430 526350
rect 543498 526294 543554 526350
rect 543622 526294 543678 526350
rect 543250 526170 543306 526226
rect 543374 526170 543430 526226
rect 543498 526170 543554 526226
rect 543622 526170 543678 526226
rect 543250 526046 543306 526102
rect 543374 526046 543430 526102
rect 543498 526046 543554 526102
rect 543622 526046 543678 526102
rect 543250 525922 543306 525978
rect 543374 525922 543430 525978
rect 543498 525922 543554 525978
rect 543622 525922 543678 525978
rect 543250 508294 543306 508350
rect 543374 508294 543430 508350
rect 543498 508294 543554 508350
rect 543622 508294 543678 508350
rect 543250 508170 543306 508226
rect 543374 508170 543430 508226
rect 543498 508170 543554 508226
rect 543622 508170 543678 508226
rect 543250 508046 543306 508102
rect 543374 508046 543430 508102
rect 543498 508046 543554 508102
rect 543622 508046 543678 508102
rect 543250 507922 543306 507978
rect 543374 507922 543430 507978
rect 543498 507922 543554 507978
rect 543622 507922 543678 507978
rect 543250 490294 543306 490350
rect 543374 490294 543430 490350
rect 543498 490294 543554 490350
rect 543622 490294 543678 490350
rect 543250 490170 543306 490226
rect 543374 490170 543430 490226
rect 543498 490170 543554 490226
rect 543622 490170 543678 490226
rect 543250 490046 543306 490102
rect 543374 490046 543430 490102
rect 543498 490046 543554 490102
rect 543622 490046 543678 490102
rect 543250 489922 543306 489978
rect 543374 489922 543430 489978
rect 543498 489922 543554 489978
rect 543622 489922 543678 489978
rect 543250 472294 543306 472350
rect 543374 472294 543430 472350
rect 543498 472294 543554 472350
rect 543622 472294 543678 472350
rect 543250 472170 543306 472226
rect 543374 472170 543430 472226
rect 543498 472170 543554 472226
rect 543622 472170 543678 472226
rect 543250 472046 543306 472102
rect 543374 472046 543430 472102
rect 543498 472046 543554 472102
rect 543622 472046 543678 472102
rect 543250 471922 543306 471978
rect 543374 471922 543430 471978
rect 543498 471922 543554 471978
rect 543622 471922 543678 471978
rect 543250 454294 543306 454350
rect 543374 454294 543430 454350
rect 543498 454294 543554 454350
rect 543622 454294 543678 454350
rect 543250 454170 543306 454226
rect 543374 454170 543430 454226
rect 543498 454170 543554 454226
rect 543622 454170 543678 454226
rect 543250 454046 543306 454102
rect 543374 454046 543430 454102
rect 543498 454046 543554 454102
rect 543622 454046 543678 454102
rect 543250 453922 543306 453978
rect 543374 453922 543430 453978
rect 543498 453922 543554 453978
rect 543622 453922 543678 453978
rect 543250 436294 543306 436350
rect 543374 436294 543430 436350
rect 543498 436294 543554 436350
rect 543622 436294 543678 436350
rect 543250 436170 543306 436226
rect 543374 436170 543430 436226
rect 543498 436170 543554 436226
rect 543622 436170 543678 436226
rect 543250 436046 543306 436102
rect 543374 436046 543430 436102
rect 543498 436046 543554 436102
rect 543622 436046 543678 436102
rect 543250 435922 543306 435978
rect 543374 435922 543430 435978
rect 543498 435922 543554 435978
rect 543622 435922 543678 435978
rect 543250 418294 543306 418350
rect 543374 418294 543430 418350
rect 543498 418294 543554 418350
rect 543622 418294 543678 418350
rect 543250 418170 543306 418226
rect 543374 418170 543430 418226
rect 543498 418170 543554 418226
rect 543622 418170 543678 418226
rect 543250 418046 543306 418102
rect 543374 418046 543430 418102
rect 543498 418046 543554 418102
rect 543622 418046 543678 418102
rect 543250 417922 543306 417978
rect 543374 417922 543430 417978
rect 543498 417922 543554 417978
rect 543622 417922 543678 417978
rect 543250 400294 543306 400350
rect 543374 400294 543430 400350
rect 543498 400294 543554 400350
rect 543622 400294 543678 400350
rect 543250 400170 543306 400226
rect 543374 400170 543430 400226
rect 543498 400170 543554 400226
rect 543622 400170 543678 400226
rect 543250 400046 543306 400102
rect 543374 400046 543430 400102
rect 543498 400046 543554 400102
rect 543622 400046 543678 400102
rect 543250 399922 543306 399978
rect 543374 399922 543430 399978
rect 543498 399922 543554 399978
rect 543622 399922 543678 399978
rect 543250 382294 543306 382350
rect 543374 382294 543430 382350
rect 543498 382294 543554 382350
rect 543622 382294 543678 382350
rect 543250 382170 543306 382226
rect 543374 382170 543430 382226
rect 543498 382170 543554 382226
rect 543622 382170 543678 382226
rect 543250 382046 543306 382102
rect 543374 382046 543430 382102
rect 543498 382046 543554 382102
rect 543622 382046 543678 382102
rect 543250 381922 543306 381978
rect 543374 381922 543430 381978
rect 543498 381922 543554 381978
rect 543622 381922 543678 381978
rect 543250 364294 543306 364350
rect 543374 364294 543430 364350
rect 543498 364294 543554 364350
rect 543622 364294 543678 364350
rect 543250 364170 543306 364226
rect 543374 364170 543430 364226
rect 543498 364170 543554 364226
rect 543622 364170 543678 364226
rect 543250 364046 543306 364102
rect 543374 364046 543430 364102
rect 543498 364046 543554 364102
rect 543622 364046 543678 364102
rect 543250 363922 543306 363978
rect 543374 363922 543430 363978
rect 543498 363922 543554 363978
rect 543622 363922 543678 363978
rect 543250 346294 543306 346350
rect 543374 346294 543430 346350
rect 543498 346294 543554 346350
rect 543622 346294 543678 346350
rect 543250 346170 543306 346226
rect 543374 346170 543430 346226
rect 543498 346170 543554 346226
rect 543622 346170 543678 346226
rect 543250 346046 543306 346102
rect 543374 346046 543430 346102
rect 543498 346046 543554 346102
rect 543622 346046 543678 346102
rect 543250 345922 543306 345978
rect 543374 345922 543430 345978
rect 543498 345922 543554 345978
rect 543622 345922 543678 345978
rect 543250 328294 543306 328350
rect 543374 328294 543430 328350
rect 543498 328294 543554 328350
rect 543622 328294 543678 328350
rect 543250 328170 543306 328226
rect 543374 328170 543430 328226
rect 543498 328170 543554 328226
rect 543622 328170 543678 328226
rect 543250 328046 543306 328102
rect 543374 328046 543430 328102
rect 543498 328046 543554 328102
rect 543622 328046 543678 328102
rect 543250 327922 543306 327978
rect 543374 327922 543430 327978
rect 543498 327922 543554 327978
rect 543622 327922 543678 327978
rect 543250 310294 543306 310350
rect 543374 310294 543430 310350
rect 543498 310294 543554 310350
rect 543622 310294 543678 310350
rect 543250 310170 543306 310226
rect 543374 310170 543430 310226
rect 543498 310170 543554 310226
rect 543622 310170 543678 310226
rect 543250 310046 543306 310102
rect 543374 310046 543430 310102
rect 543498 310046 543554 310102
rect 543622 310046 543678 310102
rect 543250 309922 543306 309978
rect 543374 309922 543430 309978
rect 543498 309922 543554 309978
rect 543622 309922 543678 309978
rect 543250 292294 543306 292350
rect 543374 292294 543430 292350
rect 543498 292294 543554 292350
rect 543622 292294 543678 292350
rect 543250 292170 543306 292226
rect 543374 292170 543430 292226
rect 543498 292170 543554 292226
rect 543622 292170 543678 292226
rect 543250 292046 543306 292102
rect 543374 292046 543430 292102
rect 543498 292046 543554 292102
rect 543622 292046 543678 292102
rect 543250 291922 543306 291978
rect 543374 291922 543430 291978
rect 543498 291922 543554 291978
rect 543622 291922 543678 291978
rect 543250 274294 543306 274350
rect 543374 274294 543430 274350
rect 543498 274294 543554 274350
rect 543622 274294 543678 274350
rect 543250 274170 543306 274226
rect 543374 274170 543430 274226
rect 543498 274170 543554 274226
rect 543622 274170 543678 274226
rect 543250 274046 543306 274102
rect 543374 274046 543430 274102
rect 543498 274046 543554 274102
rect 543622 274046 543678 274102
rect 543250 273922 543306 273978
rect 543374 273922 543430 273978
rect 543498 273922 543554 273978
rect 543622 273922 543678 273978
rect 543250 256294 543306 256350
rect 543374 256294 543430 256350
rect 543498 256294 543554 256350
rect 543622 256294 543678 256350
rect 543250 256170 543306 256226
rect 543374 256170 543430 256226
rect 543498 256170 543554 256226
rect 543622 256170 543678 256226
rect 543250 256046 543306 256102
rect 543374 256046 543430 256102
rect 543498 256046 543554 256102
rect 543622 256046 543678 256102
rect 543250 255922 543306 255978
rect 543374 255922 543430 255978
rect 543498 255922 543554 255978
rect 543622 255922 543678 255978
rect 543250 238294 543306 238350
rect 543374 238294 543430 238350
rect 543498 238294 543554 238350
rect 543622 238294 543678 238350
rect 543250 238170 543306 238226
rect 543374 238170 543430 238226
rect 543498 238170 543554 238226
rect 543622 238170 543678 238226
rect 543250 238046 543306 238102
rect 543374 238046 543430 238102
rect 543498 238046 543554 238102
rect 543622 238046 543678 238102
rect 543250 237922 543306 237978
rect 543374 237922 543430 237978
rect 543498 237922 543554 237978
rect 543622 237922 543678 237978
rect 543250 220294 543306 220350
rect 543374 220294 543430 220350
rect 543498 220294 543554 220350
rect 543622 220294 543678 220350
rect 543250 220170 543306 220226
rect 543374 220170 543430 220226
rect 543498 220170 543554 220226
rect 543622 220170 543678 220226
rect 543250 220046 543306 220102
rect 543374 220046 543430 220102
rect 543498 220046 543554 220102
rect 543622 220046 543678 220102
rect 543250 219922 543306 219978
rect 543374 219922 543430 219978
rect 543498 219922 543554 219978
rect 543622 219922 543678 219978
rect 543250 202294 543306 202350
rect 543374 202294 543430 202350
rect 543498 202294 543554 202350
rect 543622 202294 543678 202350
rect 543250 202170 543306 202226
rect 543374 202170 543430 202226
rect 543498 202170 543554 202226
rect 543622 202170 543678 202226
rect 543250 202046 543306 202102
rect 543374 202046 543430 202102
rect 543498 202046 543554 202102
rect 543622 202046 543678 202102
rect 543250 201922 543306 201978
rect 543374 201922 543430 201978
rect 543498 201922 543554 201978
rect 543622 201922 543678 201978
rect 543250 184294 543306 184350
rect 543374 184294 543430 184350
rect 543498 184294 543554 184350
rect 543622 184294 543678 184350
rect 543250 184170 543306 184226
rect 543374 184170 543430 184226
rect 543498 184170 543554 184226
rect 543622 184170 543678 184226
rect 543250 184046 543306 184102
rect 543374 184046 543430 184102
rect 543498 184046 543554 184102
rect 543622 184046 543678 184102
rect 543250 183922 543306 183978
rect 543374 183922 543430 183978
rect 543498 183922 543554 183978
rect 543622 183922 543678 183978
rect 543250 166294 543306 166350
rect 543374 166294 543430 166350
rect 543498 166294 543554 166350
rect 543622 166294 543678 166350
rect 543250 166170 543306 166226
rect 543374 166170 543430 166226
rect 543498 166170 543554 166226
rect 543622 166170 543678 166226
rect 543250 166046 543306 166102
rect 543374 166046 543430 166102
rect 543498 166046 543554 166102
rect 543622 166046 543678 166102
rect 543250 165922 543306 165978
rect 543374 165922 543430 165978
rect 543498 165922 543554 165978
rect 543622 165922 543678 165978
rect 543250 148294 543306 148350
rect 543374 148294 543430 148350
rect 543498 148294 543554 148350
rect 543622 148294 543678 148350
rect 543250 148170 543306 148226
rect 543374 148170 543430 148226
rect 543498 148170 543554 148226
rect 543622 148170 543678 148226
rect 543250 148046 543306 148102
rect 543374 148046 543430 148102
rect 543498 148046 543554 148102
rect 543622 148046 543678 148102
rect 543250 147922 543306 147978
rect 543374 147922 543430 147978
rect 543498 147922 543554 147978
rect 543622 147922 543678 147978
rect 543250 130294 543306 130350
rect 543374 130294 543430 130350
rect 543498 130294 543554 130350
rect 543622 130294 543678 130350
rect 543250 130170 543306 130226
rect 543374 130170 543430 130226
rect 543498 130170 543554 130226
rect 543622 130170 543678 130226
rect 543250 130046 543306 130102
rect 543374 130046 543430 130102
rect 543498 130046 543554 130102
rect 543622 130046 543678 130102
rect 543250 129922 543306 129978
rect 543374 129922 543430 129978
rect 543498 129922 543554 129978
rect 543622 129922 543678 129978
rect 543250 112294 543306 112350
rect 543374 112294 543430 112350
rect 543498 112294 543554 112350
rect 543622 112294 543678 112350
rect 543250 112170 543306 112226
rect 543374 112170 543430 112226
rect 543498 112170 543554 112226
rect 543622 112170 543678 112226
rect 543250 112046 543306 112102
rect 543374 112046 543430 112102
rect 543498 112046 543554 112102
rect 543622 112046 543678 112102
rect 543250 111922 543306 111978
rect 543374 111922 543430 111978
rect 543498 111922 543554 111978
rect 543622 111922 543678 111978
rect 543250 94294 543306 94350
rect 543374 94294 543430 94350
rect 543498 94294 543554 94350
rect 543622 94294 543678 94350
rect 543250 94170 543306 94226
rect 543374 94170 543430 94226
rect 543498 94170 543554 94226
rect 543622 94170 543678 94226
rect 543250 94046 543306 94102
rect 543374 94046 543430 94102
rect 543498 94046 543554 94102
rect 543622 94046 543678 94102
rect 543250 93922 543306 93978
rect 543374 93922 543430 93978
rect 543498 93922 543554 93978
rect 543622 93922 543678 93978
rect 543250 76294 543306 76350
rect 543374 76294 543430 76350
rect 543498 76294 543554 76350
rect 543622 76294 543678 76350
rect 543250 76170 543306 76226
rect 543374 76170 543430 76226
rect 543498 76170 543554 76226
rect 543622 76170 543678 76226
rect 543250 76046 543306 76102
rect 543374 76046 543430 76102
rect 543498 76046 543554 76102
rect 543622 76046 543678 76102
rect 543250 75922 543306 75978
rect 543374 75922 543430 75978
rect 543498 75922 543554 75978
rect 543622 75922 543678 75978
rect 543250 58294 543306 58350
rect 543374 58294 543430 58350
rect 543498 58294 543554 58350
rect 543622 58294 543678 58350
rect 543250 58170 543306 58226
rect 543374 58170 543430 58226
rect 543498 58170 543554 58226
rect 543622 58170 543678 58226
rect 543250 58046 543306 58102
rect 543374 58046 543430 58102
rect 543498 58046 543554 58102
rect 543622 58046 543678 58102
rect 543250 57922 543306 57978
rect 543374 57922 543430 57978
rect 543498 57922 543554 57978
rect 543622 57922 543678 57978
rect 543250 40294 543306 40350
rect 543374 40294 543430 40350
rect 543498 40294 543554 40350
rect 543622 40294 543678 40350
rect 543250 40170 543306 40226
rect 543374 40170 543430 40226
rect 543498 40170 543554 40226
rect 543622 40170 543678 40226
rect 543250 40046 543306 40102
rect 543374 40046 543430 40102
rect 543498 40046 543554 40102
rect 543622 40046 543678 40102
rect 543250 39922 543306 39978
rect 543374 39922 543430 39978
rect 543498 39922 543554 39978
rect 543622 39922 543678 39978
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 546970 514294 547026 514350
rect 547094 514294 547150 514350
rect 547218 514294 547274 514350
rect 547342 514294 547398 514350
rect 546970 514170 547026 514226
rect 547094 514170 547150 514226
rect 547218 514170 547274 514226
rect 547342 514170 547398 514226
rect 546970 514046 547026 514102
rect 547094 514046 547150 514102
rect 547218 514046 547274 514102
rect 547342 514046 547398 514102
rect 546970 513922 547026 513978
rect 547094 513922 547150 513978
rect 547218 513922 547274 513978
rect 547342 513922 547398 513978
rect 546970 496294 547026 496350
rect 547094 496294 547150 496350
rect 547218 496294 547274 496350
rect 547342 496294 547398 496350
rect 546970 496170 547026 496226
rect 547094 496170 547150 496226
rect 547218 496170 547274 496226
rect 547342 496170 547398 496226
rect 546970 496046 547026 496102
rect 547094 496046 547150 496102
rect 547218 496046 547274 496102
rect 547342 496046 547398 496102
rect 546970 495922 547026 495978
rect 547094 495922 547150 495978
rect 547218 495922 547274 495978
rect 547342 495922 547398 495978
rect 546970 478294 547026 478350
rect 547094 478294 547150 478350
rect 547218 478294 547274 478350
rect 547342 478294 547398 478350
rect 546970 478170 547026 478226
rect 547094 478170 547150 478226
rect 547218 478170 547274 478226
rect 547342 478170 547398 478226
rect 546970 478046 547026 478102
rect 547094 478046 547150 478102
rect 547218 478046 547274 478102
rect 547342 478046 547398 478102
rect 546970 477922 547026 477978
rect 547094 477922 547150 477978
rect 547218 477922 547274 477978
rect 547342 477922 547398 477978
rect 546970 460294 547026 460350
rect 547094 460294 547150 460350
rect 547218 460294 547274 460350
rect 547342 460294 547398 460350
rect 546970 460170 547026 460226
rect 547094 460170 547150 460226
rect 547218 460170 547274 460226
rect 547342 460170 547398 460226
rect 546970 460046 547026 460102
rect 547094 460046 547150 460102
rect 547218 460046 547274 460102
rect 547342 460046 547398 460102
rect 546970 459922 547026 459978
rect 547094 459922 547150 459978
rect 547218 459922 547274 459978
rect 547342 459922 547398 459978
rect 546970 442294 547026 442350
rect 547094 442294 547150 442350
rect 547218 442294 547274 442350
rect 547342 442294 547398 442350
rect 546970 442170 547026 442226
rect 547094 442170 547150 442226
rect 547218 442170 547274 442226
rect 547342 442170 547398 442226
rect 546970 442046 547026 442102
rect 547094 442046 547150 442102
rect 547218 442046 547274 442102
rect 547342 442046 547398 442102
rect 546970 441922 547026 441978
rect 547094 441922 547150 441978
rect 547218 441922 547274 441978
rect 547342 441922 547398 441978
rect 546970 424294 547026 424350
rect 547094 424294 547150 424350
rect 547218 424294 547274 424350
rect 547342 424294 547398 424350
rect 546970 424170 547026 424226
rect 547094 424170 547150 424226
rect 547218 424170 547274 424226
rect 547342 424170 547398 424226
rect 546970 424046 547026 424102
rect 547094 424046 547150 424102
rect 547218 424046 547274 424102
rect 547342 424046 547398 424102
rect 546970 423922 547026 423978
rect 547094 423922 547150 423978
rect 547218 423922 547274 423978
rect 547342 423922 547398 423978
rect 546970 406294 547026 406350
rect 547094 406294 547150 406350
rect 547218 406294 547274 406350
rect 547342 406294 547398 406350
rect 546970 406170 547026 406226
rect 547094 406170 547150 406226
rect 547218 406170 547274 406226
rect 547342 406170 547398 406226
rect 546970 406046 547026 406102
rect 547094 406046 547150 406102
rect 547218 406046 547274 406102
rect 547342 406046 547398 406102
rect 546970 405922 547026 405978
rect 547094 405922 547150 405978
rect 547218 405922 547274 405978
rect 547342 405922 547398 405978
rect 546970 388294 547026 388350
rect 547094 388294 547150 388350
rect 547218 388294 547274 388350
rect 547342 388294 547398 388350
rect 546970 388170 547026 388226
rect 547094 388170 547150 388226
rect 547218 388170 547274 388226
rect 547342 388170 547398 388226
rect 546970 388046 547026 388102
rect 547094 388046 547150 388102
rect 547218 388046 547274 388102
rect 547342 388046 547398 388102
rect 546970 387922 547026 387978
rect 547094 387922 547150 387978
rect 547218 387922 547274 387978
rect 547342 387922 547398 387978
rect 546970 370294 547026 370350
rect 547094 370294 547150 370350
rect 547218 370294 547274 370350
rect 547342 370294 547398 370350
rect 546970 370170 547026 370226
rect 547094 370170 547150 370226
rect 547218 370170 547274 370226
rect 547342 370170 547398 370226
rect 546970 370046 547026 370102
rect 547094 370046 547150 370102
rect 547218 370046 547274 370102
rect 547342 370046 547398 370102
rect 546970 369922 547026 369978
rect 547094 369922 547150 369978
rect 547218 369922 547274 369978
rect 547342 369922 547398 369978
rect 546970 352294 547026 352350
rect 547094 352294 547150 352350
rect 547218 352294 547274 352350
rect 547342 352294 547398 352350
rect 546970 352170 547026 352226
rect 547094 352170 547150 352226
rect 547218 352170 547274 352226
rect 547342 352170 547398 352226
rect 546970 352046 547026 352102
rect 547094 352046 547150 352102
rect 547218 352046 547274 352102
rect 547342 352046 547398 352102
rect 546970 351922 547026 351978
rect 547094 351922 547150 351978
rect 547218 351922 547274 351978
rect 547342 351922 547398 351978
rect 546970 334294 547026 334350
rect 547094 334294 547150 334350
rect 547218 334294 547274 334350
rect 547342 334294 547398 334350
rect 546970 334170 547026 334226
rect 547094 334170 547150 334226
rect 547218 334170 547274 334226
rect 547342 334170 547398 334226
rect 546970 334046 547026 334102
rect 547094 334046 547150 334102
rect 547218 334046 547274 334102
rect 547342 334046 547398 334102
rect 546970 333922 547026 333978
rect 547094 333922 547150 333978
rect 547218 333922 547274 333978
rect 547342 333922 547398 333978
rect 546970 316294 547026 316350
rect 547094 316294 547150 316350
rect 547218 316294 547274 316350
rect 547342 316294 547398 316350
rect 546970 316170 547026 316226
rect 547094 316170 547150 316226
rect 547218 316170 547274 316226
rect 547342 316170 547398 316226
rect 546970 316046 547026 316102
rect 547094 316046 547150 316102
rect 547218 316046 547274 316102
rect 547342 316046 547398 316102
rect 546970 315922 547026 315978
rect 547094 315922 547150 315978
rect 547218 315922 547274 315978
rect 547342 315922 547398 315978
rect 546970 298294 547026 298350
rect 547094 298294 547150 298350
rect 547218 298294 547274 298350
rect 547342 298294 547398 298350
rect 546970 298170 547026 298226
rect 547094 298170 547150 298226
rect 547218 298170 547274 298226
rect 547342 298170 547398 298226
rect 546970 298046 547026 298102
rect 547094 298046 547150 298102
rect 547218 298046 547274 298102
rect 547342 298046 547398 298102
rect 546970 297922 547026 297978
rect 547094 297922 547150 297978
rect 547218 297922 547274 297978
rect 547342 297922 547398 297978
rect 546970 280294 547026 280350
rect 547094 280294 547150 280350
rect 547218 280294 547274 280350
rect 547342 280294 547398 280350
rect 546970 280170 547026 280226
rect 547094 280170 547150 280226
rect 547218 280170 547274 280226
rect 547342 280170 547398 280226
rect 546970 280046 547026 280102
rect 547094 280046 547150 280102
rect 547218 280046 547274 280102
rect 547342 280046 547398 280102
rect 546970 279922 547026 279978
rect 547094 279922 547150 279978
rect 547218 279922 547274 279978
rect 547342 279922 547398 279978
rect 546970 262294 547026 262350
rect 547094 262294 547150 262350
rect 547218 262294 547274 262350
rect 547342 262294 547398 262350
rect 546970 262170 547026 262226
rect 547094 262170 547150 262226
rect 547218 262170 547274 262226
rect 547342 262170 547398 262226
rect 546970 262046 547026 262102
rect 547094 262046 547150 262102
rect 547218 262046 547274 262102
rect 547342 262046 547398 262102
rect 546970 261922 547026 261978
rect 547094 261922 547150 261978
rect 547218 261922 547274 261978
rect 547342 261922 547398 261978
rect 546970 244294 547026 244350
rect 547094 244294 547150 244350
rect 547218 244294 547274 244350
rect 547342 244294 547398 244350
rect 546970 244170 547026 244226
rect 547094 244170 547150 244226
rect 547218 244170 547274 244226
rect 547342 244170 547398 244226
rect 546970 244046 547026 244102
rect 547094 244046 547150 244102
rect 547218 244046 547274 244102
rect 547342 244046 547398 244102
rect 546970 243922 547026 243978
rect 547094 243922 547150 243978
rect 547218 243922 547274 243978
rect 547342 243922 547398 243978
rect 546970 226294 547026 226350
rect 547094 226294 547150 226350
rect 547218 226294 547274 226350
rect 547342 226294 547398 226350
rect 546970 226170 547026 226226
rect 547094 226170 547150 226226
rect 547218 226170 547274 226226
rect 547342 226170 547398 226226
rect 546970 226046 547026 226102
rect 547094 226046 547150 226102
rect 547218 226046 547274 226102
rect 547342 226046 547398 226102
rect 546970 225922 547026 225978
rect 547094 225922 547150 225978
rect 547218 225922 547274 225978
rect 547342 225922 547398 225978
rect 546970 208294 547026 208350
rect 547094 208294 547150 208350
rect 547218 208294 547274 208350
rect 547342 208294 547398 208350
rect 546970 208170 547026 208226
rect 547094 208170 547150 208226
rect 547218 208170 547274 208226
rect 547342 208170 547398 208226
rect 546970 208046 547026 208102
rect 547094 208046 547150 208102
rect 547218 208046 547274 208102
rect 547342 208046 547398 208102
rect 546970 207922 547026 207978
rect 547094 207922 547150 207978
rect 547218 207922 547274 207978
rect 547342 207922 547398 207978
rect 546970 190294 547026 190350
rect 547094 190294 547150 190350
rect 547218 190294 547274 190350
rect 547342 190294 547398 190350
rect 546970 190170 547026 190226
rect 547094 190170 547150 190226
rect 547218 190170 547274 190226
rect 547342 190170 547398 190226
rect 546970 190046 547026 190102
rect 547094 190046 547150 190102
rect 547218 190046 547274 190102
rect 547342 190046 547398 190102
rect 546970 189922 547026 189978
rect 547094 189922 547150 189978
rect 547218 189922 547274 189978
rect 547342 189922 547398 189978
rect 546970 172294 547026 172350
rect 547094 172294 547150 172350
rect 547218 172294 547274 172350
rect 547342 172294 547398 172350
rect 546970 172170 547026 172226
rect 547094 172170 547150 172226
rect 547218 172170 547274 172226
rect 547342 172170 547398 172226
rect 546970 172046 547026 172102
rect 547094 172046 547150 172102
rect 547218 172046 547274 172102
rect 547342 172046 547398 172102
rect 546970 171922 547026 171978
rect 547094 171922 547150 171978
rect 547218 171922 547274 171978
rect 547342 171922 547398 171978
rect 546970 154294 547026 154350
rect 547094 154294 547150 154350
rect 547218 154294 547274 154350
rect 547342 154294 547398 154350
rect 546970 154170 547026 154226
rect 547094 154170 547150 154226
rect 547218 154170 547274 154226
rect 547342 154170 547398 154226
rect 546970 154046 547026 154102
rect 547094 154046 547150 154102
rect 547218 154046 547274 154102
rect 547342 154046 547398 154102
rect 546970 153922 547026 153978
rect 547094 153922 547150 153978
rect 547218 153922 547274 153978
rect 547342 153922 547398 153978
rect 546970 136294 547026 136350
rect 547094 136294 547150 136350
rect 547218 136294 547274 136350
rect 547342 136294 547398 136350
rect 546970 136170 547026 136226
rect 547094 136170 547150 136226
rect 547218 136170 547274 136226
rect 547342 136170 547398 136226
rect 546970 136046 547026 136102
rect 547094 136046 547150 136102
rect 547218 136046 547274 136102
rect 547342 136046 547398 136102
rect 546970 135922 547026 135978
rect 547094 135922 547150 135978
rect 547218 135922 547274 135978
rect 547342 135922 547398 135978
rect 546970 118294 547026 118350
rect 547094 118294 547150 118350
rect 547218 118294 547274 118350
rect 547342 118294 547398 118350
rect 546970 118170 547026 118226
rect 547094 118170 547150 118226
rect 547218 118170 547274 118226
rect 547342 118170 547398 118226
rect 546970 118046 547026 118102
rect 547094 118046 547150 118102
rect 547218 118046 547274 118102
rect 547342 118046 547398 118102
rect 546970 117922 547026 117978
rect 547094 117922 547150 117978
rect 547218 117922 547274 117978
rect 547342 117922 547398 117978
rect 546970 100294 547026 100350
rect 547094 100294 547150 100350
rect 547218 100294 547274 100350
rect 547342 100294 547398 100350
rect 546970 100170 547026 100226
rect 547094 100170 547150 100226
rect 547218 100170 547274 100226
rect 547342 100170 547398 100226
rect 546970 100046 547026 100102
rect 547094 100046 547150 100102
rect 547218 100046 547274 100102
rect 547342 100046 547398 100102
rect 546970 99922 547026 99978
rect 547094 99922 547150 99978
rect 547218 99922 547274 99978
rect 547342 99922 547398 99978
rect 546970 82294 547026 82350
rect 547094 82294 547150 82350
rect 547218 82294 547274 82350
rect 547342 82294 547398 82350
rect 546970 82170 547026 82226
rect 547094 82170 547150 82226
rect 547218 82170 547274 82226
rect 547342 82170 547398 82226
rect 546970 82046 547026 82102
rect 547094 82046 547150 82102
rect 547218 82046 547274 82102
rect 547342 82046 547398 82102
rect 546970 81922 547026 81978
rect 547094 81922 547150 81978
rect 547218 81922 547274 81978
rect 547342 81922 547398 81978
rect 546970 64294 547026 64350
rect 547094 64294 547150 64350
rect 547218 64294 547274 64350
rect 547342 64294 547398 64350
rect 546970 64170 547026 64226
rect 547094 64170 547150 64226
rect 547218 64170 547274 64226
rect 547342 64170 547398 64226
rect 546970 64046 547026 64102
rect 547094 64046 547150 64102
rect 547218 64046 547274 64102
rect 547342 64046 547398 64102
rect 546970 63922 547026 63978
rect 547094 63922 547150 63978
rect 547218 63922 547274 63978
rect 547342 63922 547398 63978
rect 546970 46294 547026 46350
rect 547094 46294 547150 46350
rect 547218 46294 547274 46350
rect 547342 46294 547398 46350
rect 546970 46170 547026 46226
rect 547094 46170 547150 46226
rect 547218 46170 547274 46226
rect 547342 46170 547398 46226
rect 546970 46046 547026 46102
rect 547094 46046 547150 46102
rect 547218 46046 547274 46102
rect 547342 46046 547398 46102
rect 546970 45922 547026 45978
rect 547094 45922 547150 45978
rect 547218 45922 547274 45978
rect 547342 45922 547398 45978
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 561250 472294 561306 472350
rect 561374 472294 561430 472350
rect 561498 472294 561554 472350
rect 561622 472294 561678 472350
rect 561250 472170 561306 472226
rect 561374 472170 561430 472226
rect 561498 472170 561554 472226
rect 561622 472170 561678 472226
rect 561250 472046 561306 472102
rect 561374 472046 561430 472102
rect 561498 472046 561554 472102
rect 561622 472046 561678 472102
rect 561250 471922 561306 471978
rect 561374 471922 561430 471978
rect 561498 471922 561554 471978
rect 561622 471922 561678 471978
rect 561250 454294 561306 454350
rect 561374 454294 561430 454350
rect 561498 454294 561554 454350
rect 561622 454294 561678 454350
rect 561250 454170 561306 454226
rect 561374 454170 561430 454226
rect 561498 454170 561554 454226
rect 561622 454170 561678 454226
rect 561250 454046 561306 454102
rect 561374 454046 561430 454102
rect 561498 454046 561554 454102
rect 561622 454046 561678 454102
rect 561250 453922 561306 453978
rect 561374 453922 561430 453978
rect 561498 453922 561554 453978
rect 561622 453922 561678 453978
rect 561250 436294 561306 436350
rect 561374 436294 561430 436350
rect 561498 436294 561554 436350
rect 561622 436294 561678 436350
rect 561250 436170 561306 436226
rect 561374 436170 561430 436226
rect 561498 436170 561554 436226
rect 561622 436170 561678 436226
rect 561250 436046 561306 436102
rect 561374 436046 561430 436102
rect 561498 436046 561554 436102
rect 561622 436046 561678 436102
rect 561250 435922 561306 435978
rect 561374 435922 561430 435978
rect 561498 435922 561554 435978
rect 561622 435922 561678 435978
rect 561250 418294 561306 418350
rect 561374 418294 561430 418350
rect 561498 418294 561554 418350
rect 561622 418294 561678 418350
rect 561250 418170 561306 418226
rect 561374 418170 561430 418226
rect 561498 418170 561554 418226
rect 561622 418170 561678 418226
rect 561250 418046 561306 418102
rect 561374 418046 561430 418102
rect 561498 418046 561554 418102
rect 561622 418046 561678 418102
rect 561250 417922 561306 417978
rect 561374 417922 561430 417978
rect 561498 417922 561554 417978
rect 561622 417922 561678 417978
rect 561250 400294 561306 400350
rect 561374 400294 561430 400350
rect 561498 400294 561554 400350
rect 561622 400294 561678 400350
rect 561250 400170 561306 400226
rect 561374 400170 561430 400226
rect 561498 400170 561554 400226
rect 561622 400170 561678 400226
rect 561250 400046 561306 400102
rect 561374 400046 561430 400102
rect 561498 400046 561554 400102
rect 561622 400046 561678 400102
rect 561250 399922 561306 399978
rect 561374 399922 561430 399978
rect 561498 399922 561554 399978
rect 561622 399922 561678 399978
rect 561250 382294 561306 382350
rect 561374 382294 561430 382350
rect 561498 382294 561554 382350
rect 561622 382294 561678 382350
rect 561250 382170 561306 382226
rect 561374 382170 561430 382226
rect 561498 382170 561554 382226
rect 561622 382170 561678 382226
rect 561250 382046 561306 382102
rect 561374 382046 561430 382102
rect 561498 382046 561554 382102
rect 561622 382046 561678 382102
rect 561250 381922 561306 381978
rect 561374 381922 561430 381978
rect 561498 381922 561554 381978
rect 561622 381922 561678 381978
rect 561250 364294 561306 364350
rect 561374 364294 561430 364350
rect 561498 364294 561554 364350
rect 561622 364294 561678 364350
rect 561250 364170 561306 364226
rect 561374 364170 561430 364226
rect 561498 364170 561554 364226
rect 561622 364170 561678 364226
rect 561250 364046 561306 364102
rect 561374 364046 561430 364102
rect 561498 364046 561554 364102
rect 561622 364046 561678 364102
rect 561250 363922 561306 363978
rect 561374 363922 561430 363978
rect 561498 363922 561554 363978
rect 561622 363922 561678 363978
rect 561250 346294 561306 346350
rect 561374 346294 561430 346350
rect 561498 346294 561554 346350
rect 561622 346294 561678 346350
rect 561250 346170 561306 346226
rect 561374 346170 561430 346226
rect 561498 346170 561554 346226
rect 561622 346170 561678 346226
rect 561250 346046 561306 346102
rect 561374 346046 561430 346102
rect 561498 346046 561554 346102
rect 561622 346046 561678 346102
rect 561250 345922 561306 345978
rect 561374 345922 561430 345978
rect 561498 345922 561554 345978
rect 561622 345922 561678 345978
rect 561250 328294 561306 328350
rect 561374 328294 561430 328350
rect 561498 328294 561554 328350
rect 561622 328294 561678 328350
rect 561250 328170 561306 328226
rect 561374 328170 561430 328226
rect 561498 328170 561554 328226
rect 561622 328170 561678 328226
rect 561250 328046 561306 328102
rect 561374 328046 561430 328102
rect 561498 328046 561554 328102
rect 561622 328046 561678 328102
rect 561250 327922 561306 327978
rect 561374 327922 561430 327978
rect 561498 327922 561554 327978
rect 561622 327922 561678 327978
rect 561250 310294 561306 310350
rect 561374 310294 561430 310350
rect 561498 310294 561554 310350
rect 561622 310294 561678 310350
rect 561250 310170 561306 310226
rect 561374 310170 561430 310226
rect 561498 310170 561554 310226
rect 561622 310170 561678 310226
rect 561250 310046 561306 310102
rect 561374 310046 561430 310102
rect 561498 310046 561554 310102
rect 561622 310046 561678 310102
rect 561250 309922 561306 309978
rect 561374 309922 561430 309978
rect 561498 309922 561554 309978
rect 561622 309922 561678 309978
rect 561250 292294 561306 292350
rect 561374 292294 561430 292350
rect 561498 292294 561554 292350
rect 561622 292294 561678 292350
rect 561250 292170 561306 292226
rect 561374 292170 561430 292226
rect 561498 292170 561554 292226
rect 561622 292170 561678 292226
rect 561250 292046 561306 292102
rect 561374 292046 561430 292102
rect 561498 292046 561554 292102
rect 561622 292046 561678 292102
rect 561250 291922 561306 291978
rect 561374 291922 561430 291978
rect 561498 291922 561554 291978
rect 561622 291922 561678 291978
rect 561250 274294 561306 274350
rect 561374 274294 561430 274350
rect 561498 274294 561554 274350
rect 561622 274294 561678 274350
rect 561250 274170 561306 274226
rect 561374 274170 561430 274226
rect 561498 274170 561554 274226
rect 561622 274170 561678 274226
rect 561250 274046 561306 274102
rect 561374 274046 561430 274102
rect 561498 274046 561554 274102
rect 561622 274046 561678 274102
rect 561250 273922 561306 273978
rect 561374 273922 561430 273978
rect 561498 273922 561554 273978
rect 561622 273922 561678 273978
rect 561250 256294 561306 256350
rect 561374 256294 561430 256350
rect 561498 256294 561554 256350
rect 561622 256294 561678 256350
rect 561250 256170 561306 256226
rect 561374 256170 561430 256226
rect 561498 256170 561554 256226
rect 561622 256170 561678 256226
rect 561250 256046 561306 256102
rect 561374 256046 561430 256102
rect 561498 256046 561554 256102
rect 561622 256046 561678 256102
rect 561250 255922 561306 255978
rect 561374 255922 561430 255978
rect 561498 255922 561554 255978
rect 561622 255922 561678 255978
rect 561250 238294 561306 238350
rect 561374 238294 561430 238350
rect 561498 238294 561554 238350
rect 561622 238294 561678 238350
rect 561250 238170 561306 238226
rect 561374 238170 561430 238226
rect 561498 238170 561554 238226
rect 561622 238170 561678 238226
rect 561250 238046 561306 238102
rect 561374 238046 561430 238102
rect 561498 238046 561554 238102
rect 561622 238046 561678 238102
rect 561250 237922 561306 237978
rect 561374 237922 561430 237978
rect 561498 237922 561554 237978
rect 561622 237922 561678 237978
rect 561250 220294 561306 220350
rect 561374 220294 561430 220350
rect 561498 220294 561554 220350
rect 561622 220294 561678 220350
rect 561250 220170 561306 220226
rect 561374 220170 561430 220226
rect 561498 220170 561554 220226
rect 561622 220170 561678 220226
rect 561250 220046 561306 220102
rect 561374 220046 561430 220102
rect 561498 220046 561554 220102
rect 561622 220046 561678 220102
rect 561250 219922 561306 219978
rect 561374 219922 561430 219978
rect 561498 219922 561554 219978
rect 561622 219922 561678 219978
rect 561250 202294 561306 202350
rect 561374 202294 561430 202350
rect 561498 202294 561554 202350
rect 561622 202294 561678 202350
rect 561250 202170 561306 202226
rect 561374 202170 561430 202226
rect 561498 202170 561554 202226
rect 561622 202170 561678 202226
rect 561250 202046 561306 202102
rect 561374 202046 561430 202102
rect 561498 202046 561554 202102
rect 561622 202046 561678 202102
rect 561250 201922 561306 201978
rect 561374 201922 561430 201978
rect 561498 201922 561554 201978
rect 561622 201922 561678 201978
rect 561250 184294 561306 184350
rect 561374 184294 561430 184350
rect 561498 184294 561554 184350
rect 561622 184294 561678 184350
rect 561250 184170 561306 184226
rect 561374 184170 561430 184226
rect 561498 184170 561554 184226
rect 561622 184170 561678 184226
rect 561250 184046 561306 184102
rect 561374 184046 561430 184102
rect 561498 184046 561554 184102
rect 561622 184046 561678 184102
rect 561250 183922 561306 183978
rect 561374 183922 561430 183978
rect 561498 183922 561554 183978
rect 561622 183922 561678 183978
rect 561250 166294 561306 166350
rect 561374 166294 561430 166350
rect 561498 166294 561554 166350
rect 561622 166294 561678 166350
rect 561250 166170 561306 166226
rect 561374 166170 561430 166226
rect 561498 166170 561554 166226
rect 561622 166170 561678 166226
rect 561250 166046 561306 166102
rect 561374 166046 561430 166102
rect 561498 166046 561554 166102
rect 561622 166046 561678 166102
rect 561250 165922 561306 165978
rect 561374 165922 561430 165978
rect 561498 165922 561554 165978
rect 561622 165922 561678 165978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 564970 496294 565026 496350
rect 565094 496294 565150 496350
rect 565218 496294 565274 496350
rect 565342 496294 565398 496350
rect 564970 496170 565026 496226
rect 565094 496170 565150 496226
rect 565218 496170 565274 496226
rect 565342 496170 565398 496226
rect 564970 496046 565026 496102
rect 565094 496046 565150 496102
rect 565218 496046 565274 496102
rect 565342 496046 565398 496102
rect 564970 495922 565026 495978
rect 565094 495922 565150 495978
rect 565218 495922 565274 495978
rect 565342 495922 565398 495978
rect 564970 478294 565026 478350
rect 565094 478294 565150 478350
rect 565218 478294 565274 478350
rect 565342 478294 565398 478350
rect 564970 478170 565026 478226
rect 565094 478170 565150 478226
rect 565218 478170 565274 478226
rect 565342 478170 565398 478226
rect 564970 478046 565026 478102
rect 565094 478046 565150 478102
rect 565218 478046 565274 478102
rect 565342 478046 565398 478102
rect 564970 477922 565026 477978
rect 565094 477922 565150 477978
rect 565218 477922 565274 477978
rect 565342 477922 565398 477978
rect 564970 460294 565026 460350
rect 565094 460294 565150 460350
rect 565218 460294 565274 460350
rect 565342 460294 565398 460350
rect 564970 460170 565026 460226
rect 565094 460170 565150 460226
rect 565218 460170 565274 460226
rect 565342 460170 565398 460226
rect 564970 460046 565026 460102
rect 565094 460046 565150 460102
rect 565218 460046 565274 460102
rect 565342 460046 565398 460102
rect 564970 459922 565026 459978
rect 565094 459922 565150 459978
rect 565218 459922 565274 459978
rect 565342 459922 565398 459978
rect 564970 442294 565026 442350
rect 565094 442294 565150 442350
rect 565218 442294 565274 442350
rect 565342 442294 565398 442350
rect 564970 442170 565026 442226
rect 565094 442170 565150 442226
rect 565218 442170 565274 442226
rect 565342 442170 565398 442226
rect 564970 442046 565026 442102
rect 565094 442046 565150 442102
rect 565218 442046 565274 442102
rect 565342 442046 565398 442102
rect 564970 441922 565026 441978
rect 565094 441922 565150 441978
rect 565218 441922 565274 441978
rect 565342 441922 565398 441978
rect 564970 424294 565026 424350
rect 565094 424294 565150 424350
rect 565218 424294 565274 424350
rect 565342 424294 565398 424350
rect 564970 424170 565026 424226
rect 565094 424170 565150 424226
rect 565218 424170 565274 424226
rect 565342 424170 565398 424226
rect 564970 424046 565026 424102
rect 565094 424046 565150 424102
rect 565218 424046 565274 424102
rect 565342 424046 565398 424102
rect 564970 423922 565026 423978
rect 565094 423922 565150 423978
rect 565218 423922 565274 423978
rect 565342 423922 565398 423978
rect 564970 406294 565026 406350
rect 565094 406294 565150 406350
rect 565218 406294 565274 406350
rect 565342 406294 565398 406350
rect 564970 406170 565026 406226
rect 565094 406170 565150 406226
rect 565218 406170 565274 406226
rect 565342 406170 565398 406226
rect 564970 406046 565026 406102
rect 565094 406046 565150 406102
rect 565218 406046 565274 406102
rect 565342 406046 565398 406102
rect 564970 405922 565026 405978
rect 565094 405922 565150 405978
rect 565218 405922 565274 405978
rect 565342 405922 565398 405978
rect 564970 388294 565026 388350
rect 565094 388294 565150 388350
rect 565218 388294 565274 388350
rect 565342 388294 565398 388350
rect 564970 388170 565026 388226
rect 565094 388170 565150 388226
rect 565218 388170 565274 388226
rect 565342 388170 565398 388226
rect 564970 388046 565026 388102
rect 565094 388046 565150 388102
rect 565218 388046 565274 388102
rect 565342 388046 565398 388102
rect 564970 387922 565026 387978
rect 565094 387922 565150 387978
rect 565218 387922 565274 387978
rect 565342 387922 565398 387978
rect 564970 370294 565026 370350
rect 565094 370294 565150 370350
rect 565218 370294 565274 370350
rect 565342 370294 565398 370350
rect 564970 370170 565026 370226
rect 565094 370170 565150 370226
rect 565218 370170 565274 370226
rect 565342 370170 565398 370226
rect 564970 370046 565026 370102
rect 565094 370046 565150 370102
rect 565218 370046 565274 370102
rect 565342 370046 565398 370102
rect 564970 369922 565026 369978
rect 565094 369922 565150 369978
rect 565218 369922 565274 369978
rect 565342 369922 565398 369978
rect 564970 352294 565026 352350
rect 565094 352294 565150 352350
rect 565218 352294 565274 352350
rect 565342 352294 565398 352350
rect 564970 352170 565026 352226
rect 565094 352170 565150 352226
rect 565218 352170 565274 352226
rect 565342 352170 565398 352226
rect 564970 352046 565026 352102
rect 565094 352046 565150 352102
rect 565218 352046 565274 352102
rect 565342 352046 565398 352102
rect 564970 351922 565026 351978
rect 565094 351922 565150 351978
rect 565218 351922 565274 351978
rect 565342 351922 565398 351978
rect 564970 334294 565026 334350
rect 565094 334294 565150 334350
rect 565218 334294 565274 334350
rect 565342 334294 565398 334350
rect 564970 334170 565026 334226
rect 565094 334170 565150 334226
rect 565218 334170 565274 334226
rect 565342 334170 565398 334226
rect 564970 334046 565026 334102
rect 565094 334046 565150 334102
rect 565218 334046 565274 334102
rect 565342 334046 565398 334102
rect 564970 333922 565026 333978
rect 565094 333922 565150 333978
rect 565218 333922 565274 333978
rect 565342 333922 565398 333978
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298294 565026 298350
rect 565094 298294 565150 298350
rect 565218 298294 565274 298350
rect 565342 298294 565398 298350
rect 564970 298170 565026 298226
rect 565094 298170 565150 298226
rect 565218 298170 565274 298226
rect 565342 298170 565398 298226
rect 564970 298046 565026 298102
rect 565094 298046 565150 298102
rect 565218 298046 565274 298102
rect 565342 298046 565398 298102
rect 564970 297922 565026 297978
rect 565094 297922 565150 297978
rect 565218 297922 565274 297978
rect 565342 297922 565398 297978
rect 564970 280294 565026 280350
rect 565094 280294 565150 280350
rect 565218 280294 565274 280350
rect 565342 280294 565398 280350
rect 564970 280170 565026 280226
rect 565094 280170 565150 280226
rect 565218 280170 565274 280226
rect 565342 280170 565398 280226
rect 564970 280046 565026 280102
rect 565094 280046 565150 280102
rect 565218 280046 565274 280102
rect 565342 280046 565398 280102
rect 564970 279922 565026 279978
rect 565094 279922 565150 279978
rect 565218 279922 565274 279978
rect 565342 279922 565398 279978
rect 564970 262294 565026 262350
rect 565094 262294 565150 262350
rect 565218 262294 565274 262350
rect 565342 262294 565398 262350
rect 564970 262170 565026 262226
rect 565094 262170 565150 262226
rect 565218 262170 565274 262226
rect 565342 262170 565398 262226
rect 564970 262046 565026 262102
rect 565094 262046 565150 262102
rect 565218 262046 565274 262102
rect 565342 262046 565398 262102
rect 564970 261922 565026 261978
rect 565094 261922 565150 261978
rect 565218 261922 565274 261978
rect 565342 261922 565398 261978
rect 564970 244294 565026 244350
rect 565094 244294 565150 244350
rect 565218 244294 565274 244350
rect 565342 244294 565398 244350
rect 564970 244170 565026 244226
rect 565094 244170 565150 244226
rect 565218 244170 565274 244226
rect 565342 244170 565398 244226
rect 564970 244046 565026 244102
rect 565094 244046 565150 244102
rect 565218 244046 565274 244102
rect 565342 244046 565398 244102
rect 564970 243922 565026 243978
rect 565094 243922 565150 243978
rect 565218 243922 565274 243978
rect 565342 243922 565398 243978
rect 564970 226294 565026 226350
rect 565094 226294 565150 226350
rect 565218 226294 565274 226350
rect 565342 226294 565398 226350
rect 564970 226170 565026 226226
rect 565094 226170 565150 226226
rect 565218 226170 565274 226226
rect 565342 226170 565398 226226
rect 564970 226046 565026 226102
rect 565094 226046 565150 226102
rect 565218 226046 565274 226102
rect 565342 226046 565398 226102
rect 564970 225922 565026 225978
rect 565094 225922 565150 225978
rect 565218 225922 565274 225978
rect 565342 225922 565398 225978
rect 564970 208294 565026 208350
rect 565094 208294 565150 208350
rect 565218 208294 565274 208350
rect 565342 208294 565398 208350
rect 564970 208170 565026 208226
rect 565094 208170 565150 208226
rect 565218 208170 565274 208226
rect 565342 208170 565398 208226
rect 564970 208046 565026 208102
rect 565094 208046 565150 208102
rect 565218 208046 565274 208102
rect 565342 208046 565398 208102
rect 564970 207922 565026 207978
rect 565094 207922 565150 207978
rect 565218 207922 565274 207978
rect 565342 207922 565398 207978
rect 564970 190294 565026 190350
rect 565094 190294 565150 190350
rect 565218 190294 565274 190350
rect 565342 190294 565398 190350
rect 564970 190170 565026 190226
rect 565094 190170 565150 190226
rect 565218 190170 565274 190226
rect 565342 190170 565398 190226
rect 564970 190046 565026 190102
rect 565094 190046 565150 190102
rect 565218 190046 565274 190102
rect 565342 190046 565398 190102
rect 564970 189922 565026 189978
rect 565094 189922 565150 189978
rect 565218 189922 565274 189978
rect 565342 189922 565398 189978
rect 564970 172294 565026 172350
rect 565094 172294 565150 172350
rect 565218 172294 565274 172350
rect 565342 172294 565398 172350
rect 564970 172170 565026 172226
rect 565094 172170 565150 172226
rect 565218 172170 565274 172226
rect 565342 172170 565398 172226
rect 564970 172046 565026 172102
rect 565094 172046 565150 172102
rect 565218 172046 565274 172102
rect 565342 172046 565398 172102
rect 564970 171922 565026 171978
rect 565094 171922 565150 171978
rect 565218 171922 565274 171978
rect 565342 171922 565398 171978
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 579250 472294 579306 472350
rect 579374 472294 579430 472350
rect 579498 472294 579554 472350
rect 579622 472294 579678 472350
rect 579250 472170 579306 472226
rect 579374 472170 579430 472226
rect 579498 472170 579554 472226
rect 579622 472170 579678 472226
rect 579250 472046 579306 472102
rect 579374 472046 579430 472102
rect 579498 472046 579554 472102
rect 579622 472046 579678 472102
rect 579250 471922 579306 471978
rect 579374 471922 579430 471978
rect 579498 471922 579554 471978
rect 579622 471922 579678 471978
rect 579250 454294 579306 454350
rect 579374 454294 579430 454350
rect 579498 454294 579554 454350
rect 579622 454294 579678 454350
rect 579250 454170 579306 454226
rect 579374 454170 579430 454226
rect 579498 454170 579554 454226
rect 579622 454170 579678 454226
rect 579250 454046 579306 454102
rect 579374 454046 579430 454102
rect 579498 454046 579554 454102
rect 579622 454046 579678 454102
rect 579250 453922 579306 453978
rect 579374 453922 579430 453978
rect 579498 453922 579554 453978
rect 579622 453922 579678 453978
rect 579250 436294 579306 436350
rect 579374 436294 579430 436350
rect 579498 436294 579554 436350
rect 579622 436294 579678 436350
rect 579250 436170 579306 436226
rect 579374 436170 579430 436226
rect 579498 436170 579554 436226
rect 579622 436170 579678 436226
rect 579250 436046 579306 436102
rect 579374 436046 579430 436102
rect 579498 436046 579554 436102
rect 579622 436046 579678 436102
rect 579250 435922 579306 435978
rect 579374 435922 579430 435978
rect 579498 435922 579554 435978
rect 579622 435922 579678 435978
rect 579250 418294 579306 418350
rect 579374 418294 579430 418350
rect 579498 418294 579554 418350
rect 579622 418294 579678 418350
rect 579250 418170 579306 418226
rect 579374 418170 579430 418226
rect 579498 418170 579554 418226
rect 579622 418170 579678 418226
rect 579250 418046 579306 418102
rect 579374 418046 579430 418102
rect 579498 418046 579554 418102
rect 579622 418046 579678 418102
rect 579250 417922 579306 417978
rect 579374 417922 579430 417978
rect 579498 417922 579554 417978
rect 579622 417922 579678 417978
rect 579250 400294 579306 400350
rect 579374 400294 579430 400350
rect 579498 400294 579554 400350
rect 579622 400294 579678 400350
rect 579250 400170 579306 400226
rect 579374 400170 579430 400226
rect 579498 400170 579554 400226
rect 579622 400170 579678 400226
rect 579250 400046 579306 400102
rect 579374 400046 579430 400102
rect 579498 400046 579554 400102
rect 579622 400046 579678 400102
rect 579250 399922 579306 399978
rect 579374 399922 579430 399978
rect 579498 399922 579554 399978
rect 579622 399922 579678 399978
rect 579250 382294 579306 382350
rect 579374 382294 579430 382350
rect 579498 382294 579554 382350
rect 579622 382294 579678 382350
rect 579250 382170 579306 382226
rect 579374 382170 579430 382226
rect 579498 382170 579554 382226
rect 579622 382170 579678 382226
rect 579250 382046 579306 382102
rect 579374 382046 579430 382102
rect 579498 382046 579554 382102
rect 579622 382046 579678 382102
rect 579250 381922 579306 381978
rect 579374 381922 579430 381978
rect 579498 381922 579554 381978
rect 579622 381922 579678 381978
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 579250 58294 579306 58350
rect 579374 58294 579430 58350
rect 579498 58294 579554 58350
rect 579622 58294 579678 58350
rect 579250 58170 579306 58226
rect 579374 58170 579430 58226
rect 579498 58170 579554 58226
rect 579622 58170 579678 58226
rect 579250 58046 579306 58102
rect 579374 58046 579430 58102
rect 579498 58046 579554 58102
rect 579622 58046 579678 58102
rect 579250 57922 579306 57978
rect 579374 57922 579430 57978
rect 579498 57922 579554 57978
rect 579622 57922 579678 57978
rect 579250 40294 579306 40350
rect 579374 40294 579430 40350
rect 579498 40294 579554 40350
rect 579622 40294 579678 40350
rect 579250 40170 579306 40226
rect 579374 40170 579430 40226
rect 579498 40170 579554 40226
rect 579622 40170 579678 40226
rect 579250 40046 579306 40102
rect 579374 40046 579430 40102
rect 579498 40046 579554 40102
rect 579622 40046 579678 40102
rect 579250 39922 579306 39978
rect 579374 39922 579430 39978
rect 579498 39922 579554 39978
rect 579622 39922 579678 39978
rect 579250 22294 579306 22350
rect 579374 22294 579430 22350
rect 579498 22294 579554 22350
rect 579622 22294 579678 22350
rect 579250 22170 579306 22226
rect 579374 22170 579430 22226
rect 579498 22170 579554 22226
rect 579622 22170 579678 22226
rect 579250 22046 579306 22102
rect 579374 22046 579430 22102
rect 579498 22046 579554 22102
rect 579622 22046 579678 22102
rect 579250 21922 579306 21978
rect 579374 21922 579430 21978
rect 579498 21922 579554 21978
rect 579622 21922 579678 21978
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 582970 478294 583026 478350
rect 583094 478294 583150 478350
rect 583218 478294 583274 478350
rect 583342 478294 583398 478350
rect 582970 478170 583026 478226
rect 583094 478170 583150 478226
rect 583218 478170 583274 478226
rect 583342 478170 583398 478226
rect 582970 478046 583026 478102
rect 583094 478046 583150 478102
rect 583218 478046 583274 478102
rect 583342 478046 583398 478102
rect 582970 477922 583026 477978
rect 583094 477922 583150 477978
rect 583218 477922 583274 477978
rect 583342 477922 583398 477978
rect 582970 460294 583026 460350
rect 583094 460294 583150 460350
rect 583218 460294 583274 460350
rect 583342 460294 583398 460350
rect 582970 460170 583026 460226
rect 583094 460170 583150 460226
rect 583218 460170 583274 460226
rect 583342 460170 583398 460226
rect 582970 460046 583026 460102
rect 583094 460046 583150 460102
rect 583218 460046 583274 460102
rect 583342 460046 583398 460102
rect 582970 459922 583026 459978
rect 583094 459922 583150 459978
rect 583218 459922 583274 459978
rect 583342 459922 583398 459978
rect 582970 442294 583026 442350
rect 583094 442294 583150 442350
rect 583218 442294 583274 442350
rect 583342 442294 583398 442350
rect 582970 442170 583026 442226
rect 583094 442170 583150 442226
rect 583218 442170 583274 442226
rect 583342 442170 583398 442226
rect 582970 442046 583026 442102
rect 583094 442046 583150 442102
rect 583218 442046 583274 442102
rect 583342 442046 583398 442102
rect 582970 441922 583026 441978
rect 583094 441922 583150 441978
rect 583218 441922 583274 441978
rect 583342 441922 583398 441978
rect 582970 424294 583026 424350
rect 583094 424294 583150 424350
rect 583218 424294 583274 424350
rect 583342 424294 583398 424350
rect 582970 424170 583026 424226
rect 583094 424170 583150 424226
rect 583218 424170 583274 424226
rect 583342 424170 583398 424226
rect 582970 424046 583026 424102
rect 583094 424046 583150 424102
rect 583218 424046 583274 424102
rect 583342 424046 583398 424102
rect 582970 423922 583026 423978
rect 583094 423922 583150 423978
rect 583218 423922 583274 423978
rect 583342 423922 583398 423978
rect 582970 406294 583026 406350
rect 583094 406294 583150 406350
rect 583218 406294 583274 406350
rect 583342 406294 583398 406350
rect 582970 406170 583026 406226
rect 583094 406170 583150 406226
rect 583218 406170 583274 406226
rect 583342 406170 583398 406226
rect 582970 406046 583026 406102
rect 583094 406046 583150 406102
rect 583218 406046 583274 406102
rect 583342 406046 583398 406102
rect 582970 405922 583026 405978
rect 583094 405922 583150 405978
rect 583218 405922 583274 405978
rect 583342 405922 583398 405978
rect 582970 388294 583026 388350
rect 583094 388294 583150 388350
rect 583218 388294 583274 388350
rect 583342 388294 583398 388350
rect 582970 388170 583026 388226
rect 583094 388170 583150 388226
rect 583218 388170 583274 388226
rect 583342 388170 583398 388226
rect 582970 388046 583026 388102
rect 583094 388046 583150 388102
rect 583218 388046 583274 388102
rect 583342 388046 583398 388102
rect 582970 387922 583026 387978
rect 583094 387922 583150 387978
rect 583218 387922 583274 387978
rect 583342 387922 583398 387978
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 204970 496350
rect 205026 496294 205094 496350
rect 205150 496294 205218 496350
rect 205274 496294 205342 496350
rect 205398 496294 222970 496350
rect 223026 496294 223094 496350
rect 223150 496294 223218 496350
rect 223274 496294 223342 496350
rect 223398 496294 240970 496350
rect 241026 496294 241094 496350
rect 241150 496294 241218 496350
rect 241274 496294 241342 496350
rect 241398 496294 258970 496350
rect 259026 496294 259094 496350
rect 259150 496294 259218 496350
rect 259274 496294 259342 496350
rect 259398 496294 276970 496350
rect 277026 496294 277094 496350
rect 277150 496294 277218 496350
rect 277274 496294 277342 496350
rect 277398 496294 294970 496350
rect 295026 496294 295094 496350
rect 295150 496294 295218 496350
rect 295274 496294 295342 496350
rect 295398 496294 312970 496350
rect 313026 496294 313094 496350
rect 313150 496294 313218 496350
rect 313274 496294 313342 496350
rect 313398 496294 330970 496350
rect 331026 496294 331094 496350
rect 331150 496294 331218 496350
rect 331274 496294 331342 496350
rect 331398 496294 348970 496350
rect 349026 496294 349094 496350
rect 349150 496294 349218 496350
rect 349274 496294 349342 496350
rect 349398 496294 366970 496350
rect 367026 496294 367094 496350
rect 367150 496294 367218 496350
rect 367274 496294 367342 496350
rect 367398 496294 384970 496350
rect 385026 496294 385094 496350
rect 385150 496294 385218 496350
rect 385274 496294 385342 496350
rect 385398 496294 402970 496350
rect 403026 496294 403094 496350
rect 403150 496294 403218 496350
rect 403274 496294 403342 496350
rect 403398 496294 420970 496350
rect 421026 496294 421094 496350
rect 421150 496294 421218 496350
rect 421274 496294 421342 496350
rect 421398 496294 438970 496350
rect 439026 496294 439094 496350
rect 439150 496294 439218 496350
rect 439274 496294 439342 496350
rect 439398 496294 456970 496350
rect 457026 496294 457094 496350
rect 457150 496294 457218 496350
rect 457274 496294 457342 496350
rect 457398 496294 474970 496350
rect 475026 496294 475094 496350
rect 475150 496294 475218 496350
rect 475274 496294 475342 496350
rect 475398 496294 492970 496350
rect 493026 496294 493094 496350
rect 493150 496294 493218 496350
rect 493274 496294 493342 496350
rect 493398 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 204970 496226
rect 205026 496170 205094 496226
rect 205150 496170 205218 496226
rect 205274 496170 205342 496226
rect 205398 496170 222970 496226
rect 223026 496170 223094 496226
rect 223150 496170 223218 496226
rect 223274 496170 223342 496226
rect 223398 496170 240970 496226
rect 241026 496170 241094 496226
rect 241150 496170 241218 496226
rect 241274 496170 241342 496226
rect 241398 496170 258970 496226
rect 259026 496170 259094 496226
rect 259150 496170 259218 496226
rect 259274 496170 259342 496226
rect 259398 496170 276970 496226
rect 277026 496170 277094 496226
rect 277150 496170 277218 496226
rect 277274 496170 277342 496226
rect 277398 496170 294970 496226
rect 295026 496170 295094 496226
rect 295150 496170 295218 496226
rect 295274 496170 295342 496226
rect 295398 496170 312970 496226
rect 313026 496170 313094 496226
rect 313150 496170 313218 496226
rect 313274 496170 313342 496226
rect 313398 496170 330970 496226
rect 331026 496170 331094 496226
rect 331150 496170 331218 496226
rect 331274 496170 331342 496226
rect 331398 496170 348970 496226
rect 349026 496170 349094 496226
rect 349150 496170 349218 496226
rect 349274 496170 349342 496226
rect 349398 496170 366970 496226
rect 367026 496170 367094 496226
rect 367150 496170 367218 496226
rect 367274 496170 367342 496226
rect 367398 496170 384970 496226
rect 385026 496170 385094 496226
rect 385150 496170 385218 496226
rect 385274 496170 385342 496226
rect 385398 496170 402970 496226
rect 403026 496170 403094 496226
rect 403150 496170 403218 496226
rect 403274 496170 403342 496226
rect 403398 496170 420970 496226
rect 421026 496170 421094 496226
rect 421150 496170 421218 496226
rect 421274 496170 421342 496226
rect 421398 496170 438970 496226
rect 439026 496170 439094 496226
rect 439150 496170 439218 496226
rect 439274 496170 439342 496226
rect 439398 496170 456970 496226
rect 457026 496170 457094 496226
rect 457150 496170 457218 496226
rect 457274 496170 457342 496226
rect 457398 496170 474970 496226
rect 475026 496170 475094 496226
rect 475150 496170 475218 496226
rect 475274 496170 475342 496226
rect 475398 496170 492970 496226
rect 493026 496170 493094 496226
rect 493150 496170 493218 496226
rect 493274 496170 493342 496226
rect 493398 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 204970 496102
rect 205026 496046 205094 496102
rect 205150 496046 205218 496102
rect 205274 496046 205342 496102
rect 205398 496046 222970 496102
rect 223026 496046 223094 496102
rect 223150 496046 223218 496102
rect 223274 496046 223342 496102
rect 223398 496046 240970 496102
rect 241026 496046 241094 496102
rect 241150 496046 241218 496102
rect 241274 496046 241342 496102
rect 241398 496046 258970 496102
rect 259026 496046 259094 496102
rect 259150 496046 259218 496102
rect 259274 496046 259342 496102
rect 259398 496046 276970 496102
rect 277026 496046 277094 496102
rect 277150 496046 277218 496102
rect 277274 496046 277342 496102
rect 277398 496046 294970 496102
rect 295026 496046 295094 496102
rect 295150 496046 295218 496102
rect 295274 496046 295342 496102
rect 295398 496046 312970 496102
rect 313026 496046 313094 496102
rect 313150 496046 313218 496102
rect 313274 496046 313342 496102
rect 313398 496046 330970 496102
rect 331026 496046 331094 496102
rect 331150 496046 331218 496102
rect 331274 496046 331342 496102
rect 331398 496046 348970 496102
rect 349026 496046 349094 496102
rect 349150 496046 349218 496102
rect 349274 496046 349342 496102
rect 349398 496046 366970 496102
rect 367026 496046 367094 496102
rect 367150 496046 367218 496102
rect 367274 496046 367342 496102
rect 367398 496046 384970 496102
rect 385026 496046 385094 496102
rect 385150 496046 385218 496102
rect 385274 496046 385342 496102
rect 385398 496046 402970 496102
rect 403026 496046 403094 496102
rect 403150 496046 403218 496102
rect 403274 496046 403342 496102
rect 403398 496046 420970 496102
rect 421026 496046 421094 496102
rect 421150 496046 421218 496102
rect 421274 496046 421342 496102
rect 421398 496046 438970 496102
rect 439026 496046 439094 496102
rect 439150 496046 439218 496102
rect 439274 496046 439342 496102
rect 439398 496046 456970 496102
rect 457026 496046 457094 496102
rect 457150 496046 457218 496102
rect 457274 496046 457342 496102
rect 457398 496046 474970 496102
rect 475026 496046 475094 496102
rect 475150 496046 475218 496102
rect 475274 496046 475342 496102
rect 475398 496046 492970 496102
rect 493026 496046 493094 496102
rect 493150 496046 493218 496102
rect 493274 496046 493342 496102
rect 493398 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 204970 495978
rect 205026 495922 205094 495978
rect 205150 495922 205218 495978
rect 205274 495922 205342 495978
rect 205398 495922 222970 495978
rect 223026 495922 223094 495978
rect 223150 495922 223218 495978
rect 223274 495922 223342 495978
rect 223398 495922 240970 495978
rect 241026 495922 241094 495978
rect 241150 495922 241218 495978
rect 241274 495922 241342 495978
rect 241398 495922 258970 495978
rect 259026 495922 259094 495978
rect 259150 495922 259218 495978
rect 259274 495922 259342 495978
rect 259398 495922 276970 495978
rect 277026 495922 277094 495978
rect 277150 495922 277218 495978
rect 277274 495922 277342 495978
rect 277398 495922 294970 495978
rect 295026 495922 295094 495978
rect 295150 495922 295218 495978
rect 295274 495922 295342 495978
rect 295398 495922 312970 495978
rect 313026 495922 313094 495978
rect 313150 495922 313218 495978
rect 313274 495922 313342 495978
rect 313398 495922 330970 495978
rect 331026 495922 331094 495978
rect 331150 495922 331218 495978
rect 331274 495922 331342 495978
rect 331398 495922 348970 495978
rect 349026 495922 349094 495978
rect 349150 495922 349218 495978
rect 349274 495922 349342 495978
rect 349398 495922 366970 495978
rect 367026 495922 367094 495978
rect 367150 495922 367218 495978
rect 367274 495922 367342 495978
rect 367398 495922 384970 495978
rect 385026 495922 385094 495978
rect 385150 495922 385218 495978
rect 385274 495922 385342 495978
rect 385398 495922 402970 495978
rect 403026 495922 403094 495978
rect 403150 495922 403218 495978
rect 403274 495922 403342 495978
rect 403398 495922 420970 495978
rect 421026 495922 421094 495978
rect 421150 495922 421218 495978
rect 421274 495922 421342 495978
rect 421398 495922 438970 495978
rect 439026 495922 439094 495978
rect 439150 495922 439218 495978
rect 439274 495922 439342 495978
rect 439398 495922 456970 495978
rect 457026 495922 457094 495978
rect 457150 495922 457218 495978
rect 457274 495922 457342 495978
rect 457398 495922 474970 495978
rect 475026 495922 475094 495978
rect 475150 495922 475218 495978
rect 475274 495922 475342 495978
rect 475398 495922 492970 495978
rect 493026 495922 493094 495978
rect 493150 495922 493218 495978
rect 493274 495922 493342 495978
rect 493398 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 219250 490350
rect 219306 490294 219374 490350
rect 219430 490294 219498 490350
rect 219554 490294 219622 490350
rect 219678 490294 237250 490350
rect 237306 490294 237374 490350
rect 237430 490294 237498 490350
rect 237554 490294 237622 490350
rect 237678 490294 255250 490350
rect 255306 490294 255374 490350
rect 255430 490294 255498 490350
rect 255554 490294 255622 490350
rect 255678 490294 273250 490350
rect 273306 490294 273374 490350
rect 273430 490294 273498 490350
rect 273554 490294 273622 490350
rect 273678 490294 291250 490350
rect 291306 490294 291374 490350
rect 291430 490294 291498 490350
rect 291554 490294 291622 490350
rect 291678 490294 309250 490350
rect 309306 490294 309374 490350
rect 309430 490294 309498 490350
rect 309554 490294 309622 490350
rect 309678 490294 327250 490350
rect 327306 490294 327374 490350
rect 327430 490294 327498 490350
rect 327554 490294 327622 490350
rect 327678 490294 345250 490350
rect 345306 490294 345374 490350
rect 345430 490294 345498 490350
rect 345554 490294 345622 490350
rect 345678 490294 363250 490350
rect 363306 490294 363374 490350
rect 363430 490294 363498 490350
rect 363554 490294 363622 490350
rect 363678 490294 381250 490350
rect 381306 490294 381374 490350
rect 381430 490294 381498 490350
rect 381554 490294 381622 490350
rect 381678 490294 399250 490350
rect 399306 490294 399374 490350
rect 399430 490294 399498 490350
rect 399554 490294 399622 490350
rect 399678 490294 417250 490350
rect 417306 490294 417374 490350
rect 417430 490294 417498 490350
rect 417554 490294 417622 490350
rect 417678 490294 435250 490350
rect 435306 490294 435374 490350
rect 435430 490294 435498 490350
rect 435554 490294 435622 490350
rect 435678 490294 453250 490350
rect 453306 490294 453374 490350
rect 453430 490294 453498 490350
rect 453554 490294 453622 490350
rect 453678 490294 471250 490350
rect 471306 490294 471374 490350
rect 471430 490294 471498 490350
rect 471554 490294 471622 490350
rect 471678 490294 489250 490350
rect 489306 490294 489374 490350
rect 489430 490294 489498 490350
rect 489554 490294 489622 490350
rect 489678 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 219250 490226
rect 219306 490170 219374 490226
rect 219430 490170 219498 490226
rect 219554 490170 219622 490226
rect 219678 490170 237250 490226
rect 237306 490170 237374 490226
rect 237430 490170 237498 490226
rect 237554 490170 237622 490226
rect 237678 490170 255250 490226
rect 255306 490170 255374 490226
rect 255430 490170 255498 490226
rect 255554 490170 255622 490226
rect 255678 490170 273250 490226
rect 273306 490170 273374 490226
rect 273430 490170 273498 490226
rect 273554 490170 273622 490226
rect 273678 490170 291250 490226
rect 291306 490170 291374 490226
rect 291430 490170 291498 490226
rect 291554 490170 291622 490226
rect 291678 490170 309250 490226
rect 309306 490170 309374 490226
rect 309430 490170 309498 490226
rect 309554 490170 309622 490226
rect 309678 490170 327250 490226
rect 327306 490170 327374 490226
rect 327430 490170 327498 490226
rect 327554 490170 327622 490226
rect 327678 490170 345250 490226
rect 345306 490170 345374 490226
rect 345430 490170 345498 490226
rect 345554 490170 345622 490226
rect 345678 490170 363250 490226
rect 363306 490170 363374 490226
rect 363430 490170 363498 490226
rect 363554 490170 363622 490226
rect 363678 490170 381250 490226
rect 381306 490170 381374 490226
rect 381430 490170 381498 490226
rect 381554 490170 381622 490226
rect 381678 490170 399250 490226
rect 399306 490170 399374 490226
rect 399430 490170 399498 490226
rect 399554 490170 399622 490226
rect 399678 490170 417250 490226
rect 417306 490170 417374 490226
rect 417430 490170 417498 490226
rect 417554 490170 417622 490226
rect 417678 490170 435250 490226
rect 435306 490170 435374 490226
rect 435430 490170 435498 490226
rect 435554 490170 435622 490226
rect 435678 490170 453250 490226
rect 453306 490170 453374 490226
rect 453430 490170 453498 490226
rect 453554 490170 453622 490226
rect 453678 490170 471250 490226
rect 471306 490170 471374 490226
rect 471430 490170 471498 490226
rect 471554 490170 471622 490226
rect 471678 490170 489250 490226
rect 489306 490170 489374 490226
rect 489430 490170 489498 490226
rect 489554 490170 489622 490226
rect 489678 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 219250 490102
rect 219306 490046 219374 490102
rect 219430 490046 219498 490102
rect 219554 490046 219622 490102
rect 219678 490046 237250 490102
rect 237306 490046 237374 490102
rect 237430 490046 237498 490102
rect 237554 490046 237622 490102
rect 237678 490046 255250 490102
rect 255306 490046 255374 490102
rect 255430 490046 255498 490102
rect 255554 490046 255622 490102
rect 255678 490046 273250 490102
rect 273306 490046 273374 490102
rect 273430 490046 273498 490102
rect 273554 490046 273622 490102
rect 273678 490046 291250 490102
rect 291306 490046 291374 490102
rect 291430 490046 291498 490102
rect 291554 490046 291622 490102
rect 291678 490046 309250 490102
rect 309306 490046 309374 490102
rect 309430 490046 309498 490102
rect 309554 490046 309622 490102
rect 309678 490046 327250 490102
rect 327306 490046 327374 490102
rect 327430 490046 327498 490102
rect 327554 490046 327622 490102
rect 327678 490046 345250 490102
rect 345306 490046 345374 490102
rect 345430 490046 345498 490102
rect 345554 490046 345622 490102
rect 345678 490046 363250 490102
rect 363306 490046 363374 490102
rect 363430 490046 363498 490102
rect 363554 490046 363622 490102
rect 363678 490046 381250 490102
rect 381306 490046 381374 490102
rect 381430 490046 381498 490102
rect 381554 490046 381622 490102
rect 381678 490046 399250 490102
rect 399306 490046 399374 490102
rect 399430 490046 399498 490102
rect 399554 490046 399622 490102
rect 399678 490046 417250 490102
rect 417306 490046 417374 490102
rect 417430 490046 417498 490102
rect 417554 490046 417622 490102
rect 417678 490046 435250 490102
rect 435306 490046 435374 490102
rect 435430 490046 435498 490102
rect 435554 490046 435622 490102
rect 435678 490046 453250 490102
rect 453306 490046 453374 490102
rect 453430 490046 453498 490102
rect 453554 490046 453622 490102
rect 453678 490046 471250 490102
rect 471306 490046 471374 490102
rect 471430 490046 471498 490102
rect 471554 490046 471622 490102
rect 471678 490046 489250 490102
rect 489306 490046 489374 490102
rect 489430 490046 489498 490102
rect 489554 490046 489622 490102
rect 489678 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 219250 489978
rect 219306 489922 219374 489978
rect 219430 489922 219498 489978
rect 219554 489922 219622 489978
rect 219678 489922 237250 489978
rect 237306 489922 237374 489978
rect 237430 489922 237498 489978
rect 237554 489922 237622 489978
rect 237678 489922 255250 489978
rect 255306 489922 255374 489978
rect 255430 489922 255498 489978
rect 255554 489922 255622 489978
rect 255678 489922 273250 489978
rect 273306 489922 273374 489978
rect 273430 489922 273498 489978
rect 273554 489922 273622 489978
rect 273678 489922 291250 489978
rect 291306 489922 291374 489978
rect 291430 489922 291498 489978
rect 291554 489922 291622 489978
rect 291678 489922 309250 489978
rect 309306 489922 309374 489978
rect 309430 489922 309498 489978
rect 309554 489922 309622 489978
rect 309678 489922 327250 489978
rect 327306 489922 327374 489978
rect 327430 489922 327498 489978
rect 327554 489922 327622 489978
rect 327678 489922 345250 489978
rect 345306 489922 345374 489978
rect 345430 489922 345498 489978
rect 345554 489922 345622 489978
rect 345678 489922 363250 489978
rect 363306 489922 363374 489978
rect 363430 489922 363498 489978
rect 363554 489922 363622 489978
rect 363678 489922 381250 489978
rect 381306 489922 381374 489978
rect 381430 489922 381498 489978
rect 381554 489922 381622 489978
rect 381678 489922 399250 489978
rect 399306 489922 399374 489978
rect 399430 489922 399498 489978
rect 399554 489922 399622 489978
rect 399678 489922 417250 489978
rect 417306 489922 417374 489978
rect 417430 489922 417498 489978
rect 417554 489922 417622 489978
rect 417678 489922 435250 489978
rect 435306 489922 435374 489978
rect 435430 489922 435498 489978
rect 435554 489922 435622 489978
rect 435678 489922 453250 489978
rect 453306 489922 453374 489978
rect 453430 489922 453498 489978
rect 453554 489922 453622 489978
rect 453678 489922 471250 489978
rect 471306 489922 471374 489978
rect 471430 489922 471498 489978
rect 471554 489922 471622 489978
rect 471678 489922 489250 489978
rect 489306 489922 489374 489978
rect 489430 489922 489498 489978
rect 489554 489922 489622 489978
rect 489678 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 204970 478350
rect 205026 478294 205094 478350
rect 205150 478294 205218 478350
rect 205274 478294 205342 478350
rect 205398 478294 222970 478350
rect 223026 478294 223094 478350
rect 223150 478294 223218 478350
rect 223274 478294 223342 478350
rect 223398 478294 240970 478350
rect 241026 478294 241094 478350
rect 241150 478294 241218 478350
rect 241274 478294 241342 478350
rect 241398 478294 258970 478350
rect 259026 478294 259094 478350
rect 259150 478294 259218 478350
rect 259274 478294 259342 478350
rect 259398 478294 276970 478350
rect 277026 478294 277094 478350
rect 277150 478294 277218 478350
rect 277274 478294 277342 478350
rect 277398 478294 294970 478350
rect 295026 478294 295094 478350
rect 295150 478294 295218 478350
rect 295274 478294 295342 478350
rect 295398 478294 312970 478350
rect 313026 478294 313094 478350
rect 313150 478294 313218 478350
rect 313274 478294 313342 478350
rect 313398 478294 330970 478350
rect 331026 478294 331094 478350
rect 331150 478294 331218 478350
rect 331274 478294 331342 478350
rect 331398 478294 348970 478350
rect 349026 478294 349094 478350
rect 349150 478294 349218 478350
rect 349274 478294 349342 478350
rect 349398 478294 366970 478350
rect 367026 478294 367094 478350
rect 367150 478294 367218 478350
rect 367274 478294 367342 478350
rect 367398 478294 384970 478350
rect 385026 478294 385094 478350
rect 385150 478294 385218 478350
rect 385274 478294 385342 478350
rect 385398 478294 402970 478350
rect 403026 478294 403094 478350
rect 403150 478294 403218 478350
rect 403274 478294 403342 478350
rect 403398 478294 420970 478350
rect 421026 478294 421094 478350
rect 421150 478294 421218 478350
rect 421274 478294 421342 478350
rect 421398 478294 438970 478350
rect 439026 478294 439094 478350
rect 439150 478294 439218 478350
rect 439274 478294 439342 478350
rect 439398 478294 456970 478350
rect 457026 478294 457094 478350
rect 457150 478294 457218 478350
rect 457274 478294 457342 478350
rect 457398 478294 474970 478350
rect 475026 478294 475094 478350
rect 475150 478294 475218 478350
rect 475274 478294 475342 478350
rect 475398 478294 492970 478350
rect 493026 478294 493094 478350
rect 493150 478294 493218 478350
rect 493274 478294 493342 478350
rect 493398 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 204970 478226
rect 205026 478170 205094 478226
rect 205150 478170 205218 478226
rect 205274 478170 205342 478226
rect 205398 478170 222970 478226
rect 223026 478170 223094 478226
rect 223150 478170 223218 478226
rect 223274 478170 223342 478226
rect 223398 478170 240970 478226
rect 241026 478170 241094 478226
rect 241150 478170 241218 478226
rect 241274 478170 241342 478226
rect 241398 478170 258970 478226
rect 259026 478170 259094 478226
rect 259150 478170 259218 478226
rect 259274 478170 259342 478226
rect 259398 478170 276970 478226
rect 277026 478170 277094 478226
rect 277150 478170 277218 478226
rect 277274 478170 277342 478226
rect 277398 478170 294970 478226
rect 295026 478170 295094 478226
rect 295150 478170 295218 478226
rect 295274 478170 295342 478226
rect 295398 478170 312970 478226
rect 313026 478170 313094 478226
rect 313150 478170 313218 478226
rect 313274 478170 313342 478226
rect 313398 478170 330970 478226
rect 331026 478170 331094 478226
rect 331150 478170 331218 478226
rect 331274 478170 331342 478226
rect 331398 478170 348970 478226
rect 349026 478170 349094 478226
rect 349150 478170 349218 478226
rect 349274 478170 349342 478226
rect 349398 478170 366970 478226
rect 367026 478170 367094 478226
rect 367150 478170 367218 478226
rect 367274 478170 367342 478226
rect 367398 478170 384970 478226
rect 385026 478170 385094 478226
rect 385150 478170 385218 478226
rect 385274 478170 385342 478226
rect 385398 478170 402970 478226
rect 403026 478170 403094 478226
rect 403150 478170 403218 478226
rect 403274 478170 403342 478226
rect 403398 478170 420970 478226
rect 421026 478170 421094 478226
rect 421150 478170 421218 478226
rect 421274 478170 421342 478226
rect 421398 478170 438970 478226
rect 439026 478170 439094 478226
rect 439150 478170 439218 478226
rect 439274 478170 439342 478226
rect 439398 478170 456970 478226
rect 457026 478170 457094 478226
rect 457150 478170 457218 478226
rect 457274 478170 457342 478226
rect 457398 478170 474970 478226
rect 475026 478170 475094 478226
rect 475150 478170 475218 478226
rect 475274 478170 475342 478226
rect 475398 478170 492970 478226
rect 493026 478170 493094 478226
rect 493150 478170 493218 478226
rect 493274 478170 493342 478226
rect 493398 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 204970 478102
rect 205026 478046 205094 478102
rect 205150 478046 205218 478102
rect 205274 478046 205342 478102
rect 205398 478046 222970 478102
rect 223026 478046 223094 478102
rect 223150 478046 223218 478102
rect 223274 478046 223342 478102
rect 223398 478046 240970 478102
rect 241026 478046 241094 478102
rect 241150 478046 241218 478102
rect 241274 478046 241342 478102
rect 241398 478046 258970 478102
rect 259026 478046 259094 478102
rect 259150 478046 259218 478102
rect 259274 478046 259342 478102
rect 259398 478046 276970 478102
rect 277026 478046 277094 478102
rect 277150 478046 277218 478102
rect 277274 478046 277342 478102
rect 277398 478046 294970 478102
rect 295026 478046 295094 478102
rect 295150 478046 295218 478102
rect 295274 478046 295342 478102
rect 295398 478046 312970 478102
rect 313026 478046 313094 478102
rect 313150 478046 313218 478102
rect 313274 478046 313342 478102
rect 313398 478046 330970 478102
rect 331026 478046 331094 478102
rect 331150 478046 331218 478102
rect 331274 478046 331342 478102
rect 331398 478046 348970 478102
rect 349026 478046 349094 478102
rect 349150 478046 349218 478102
rect 349274 478046 349342 478102
rect 349398 478046 366970 478102
rect 367026 478046 367094 478102
rect 367150 478046 367218 478102
rect 367274 478046 367342 478102
rect 367398 478046 384970 478102
rect 385026 478046 385094 478102
rect 385150 478046 385218 478102
rect 385274 478046 385342 478102
rect 385398 478046 402970 478102
rect 403026 478046 403094 478102
rect 403150 478046 403218 478102
rect 403274 478046 403342 478102
rect 403398 478046 420970 478102
rect 421026 478046 421094 478102
rect 421150 478046 421218 478102
rect 421274 478046 421342 478102
rect 421398 478046 438970 478102
rect 439026 478046 439094 478102
rect 439150 478046 439218 478102
rect 439274 478046 439342 478102
rect 439398 478046 456970 478102
rect 457026 478046 457094 478102
rect 457150 478046 457218 478102
rect 457274 478046 457342 478102
rect 457398 478046 474970 478102
rect 475026 478046 475094 478102
rect 475150 478046 475218 478102
rect 475274 478046 475342 478102
rect 475398 478046 492970 478102
rect 493026 478046 493094 478102
rect 493150 478046 493218 478102
rect 493274 478046 493342 478102
rect 493398 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 204970 477978
rect 205026 477922 205094 477978
rect 205150 477922 205218 477978
rect 205274 477922 205342 477978
rect 205398 477922 222970 477978
rect 223026 477922 223094 477978
rect 223150 477922 223218 477978
rect 223274 477922 223342 477978
rect 223398 477922 240970 477978
rect 241026 477922 241094 477978
rect 241150 477922 241218 477978
rect 241274 477922 241342 477978
rect 241398 477922 258970 477978
rect 259026 477922 259094 477978
rect 259150 477922 259218 477978
rect 259274 477922 259342 477978
rect 259398 477922 276970 477978
rect 277026 477922 277094 477978
rect 277150 477922 277218 477978
rect 277274 477922 277342 477978
rect 277398 477922 294970 477978
rect 295026 477922 295094 477978
rect 295150 477922 295218 477978
rect 295274 477922 295342 477978
rect 295398 477922 312970 477978
rect 313026 477922 313094 477978
rect 313150 477922 313218 477978
rect 313274 477922 313342 477978
rect 313398 477922 330970 477978
rect 331026 477922 331094 477978
rect 331150 477922 331218 477978
rect 331274 477922 331342 477978
rect 331398 477922 348970 477978
rect 349026 477922 349094 477978
rect 349150 477922 349218 477978
rect 349274 477922 349342 477978
rect 349398 477922 366970 477978
rect 367026 477922 367094 477978
rect 367150 477922 367218 477978
rect 367274 477922 367342 477978
rect 367398 477922 384970 477978
rect 385026 477922 385094 477978
rect 385150 477922 385218 477978
rect 385274 477922 385342 477978
rect 385398 477922 402970 477978
rect 403026 477922 403094 477978
rect 403150 477922 403218 477978
rect 403274 477922 403342 477978
rect 403398 477922 420970 477978
rect 421026 477922 421094 477978
rect 421150 477922 421218 477978
rect 421274 477922 421342 477978
rect 421398 477922 438970 477978
rect 439026 477922 439094 477978
rect 439150 477922 439218 477978
rect 439274 477922 439342 477978
rect 439398 477922 456970 477978
rect 457026 477922 457094 477978
rect 457150 477922 457218 477978
rect 457274 477922 457342 477978
rect 457398 477922 474970 477978
rect 475026 477922 475094 477978
rect 475150 477922 475218 477978
rect 475274 477922 475342 477978
rect 475398 477922 492970 477978
rect 493026 477922 493094 477978
rect 493150 477922 493218 477978
rect 493274 477922 493342 477978
rect 493398 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 219250 472350
rect 219306 472294 219374 472350
rect 219430 472294 219498 472350
rect 219554 472294 219622 472350
rect 219678 472294 237250 472350
rect 237306 472294 237374 472350
rect 237430 472294 237498 472350
rect 237554 472294 237622 472350
rect 237678 472294 255250 472350
rect 255306 472294 255374 472350
rect 255430 472294 255498 472350
rect 255554 472294 255622 472350
rect 255678 472294 273250 472350
rect 273306 472294 273374 472350
rect 273430 472294 273498 472350
rect 273554 472294 273622 472350
rect 273678 472294 291250 472350
rect 291306 472294 291374 472350
rect 291430 472294 291498 472350
rect 291554 472294 291622 472350
rect 291678 472294 309250 472350
rect 309306 472294 309374 472350
rect 309430 472294 309498 472350
rect 309554 472294 309622 472350
rect 309678 472294 327250 472350
rect 327306 472294 327374 472350
rect 327430 472294 327498 472350
rect 327554 472294 327622 472350
rect 327678 472294 345250 472350
rect 345306 472294 345374 472350
rect 345430 472294 345498 472350
rect 345554 472294 345622 472350
rect 345678 472294 363250 472350
rect 363306 472294 363374 472350
rect 363430 472294 363498 472350
rect 363554 472294 363622 472350
rect 363678 472294 381250 472350
rect 381306 472294 381374 472350
rect 381430 472294 381498 472350
rect 381554 472294 381622 472350
rect 381678 472294 399250 472350
rect 399306 472294 399374 472350
rect 399430 472294 399498 472350
rect 399554 472294 399622 472350
rect 399678 472294 417250 472350
rect 417306 472294 417374 472350
rect 417430 472294 417498 472350
rect 417554 472294 417622 472350
rect 417678 472294 435250 472350
rect 435306 472294 435374 472350
rect 435430 472294 435498 472350
rect 435554 472294 435622 472350
rect 435678 472294 453250 472350
rect 453306 472294 453374 472350
rect 453430 472294 453498 472350
rect 453554 472294 453622 472350
rect 453678 472294 471250 472350
rect 471306 472294 471374 472350
rect 471430 472294 471498 472350
rect 471554 472294 471622 472350
rect 471678 472294 489250 472350
rect 489306 472294 489374 472350
rect 489430 472294 489498 472350
rect 489554 472294 489622 472350
rect 489678 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 219250 472226
rect 219306 472170 219374 472226
rect 219430 472170 219498 472226
rect 219554 472170 219622 472226
rect 219678 472170 237250 472226
rect 237306 472170 237374 472226
rect 237430 472170 237498 472226
rect 237554 472170 237622 472226
rect 237678 472170 255250 472226
rect 255306 472170 255374 472226
rect 255430 472170 255498 472226
rect 255554 472170 255622 472226
rect 255678 472170 273250 472226
rect 273306 472170 273374 472226
rect 273430 472170 273498 472226
rect 273554 472170 273622 472226
rect 273678 472170 291250 472226
rect 291306 472170 291374 472226
rect 291430 472170 291498 472226
rect 291554 472170 291622 472226
rect 291678 472170 309250 472226
rect 309306 472170 309374 472226
rect 309430 472170 309498 472226
rect 309554 472170 309622 472226
rect 309678 472170 327250 472226
rect 327306 472170 327374 472226
rect 327430 472170 327498 472226
rect 327554 472170 327622 472226
rect 327678 472170 345250 472226
rect 345306 472170 345374 472226
rect 345430 472170 345498 472226
rect 345554 472170 345622 472226
rect 345678 472170 363250 472226
rect 363306 472170 363374 472226
rect 363430 472170 363498 472226
rect 363554 472170 363622 472226
rect 363678 472170 381250 472226
rect 381306 472170 381374 472226
rect 381430 472170 381498 472226
rect 381554 472170 381622 472226
rect 381678 472170 399250 472226
rect 399306 472170 399374 472226
rect 399430 472170 399498 472226
rect 399554 472170 399622 472226
rect 399678 472170 417250 472226
rect 417306 472170 417374 472226
rect 417430 472170 417498 472226
rect 417554 472170 417622 472226
rect 417678 472170 435250 472226
rect 435306 472170 435374 472226
rect 435430 472170 435498 472226
rect 435554 472170 435622 472226
rect 435678 472170 453250 472226
rect 453306 472170 453374 472226
rect 453430 472170 453498 472226
rect 453554 472170 453622 472226
rect 453678 472170 471250 472226
rect 471306 472170 471374 472226
rect 471430 472170 471498 472226
rect 471554 472170 471622 472226
rect 471678 472170 489250 472226
rect 489306 472170 489374 472226
rect 489430 472170 489498 472226
rect 489554 472170 489622 472226
rect 489678 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 219250 472102
rect 219306 472046 219374 472102
rect 219430 472046 219498 472102
rect 219554 472046 219622 472102
rect 219678 472046 237250 472102
rect 237306 472046 237374 472102
rect 237430 472046 237498 472102
rect 237554 472046 237622 472102
rect 237678 472046 255250 472102
rect 255306 472046 255374 472102
rect 255430 472046 255498 472102
rect 255554 472046 255622 472102
rect 255678 472046 273250 472102
rect 273306 472046 273374 472102
rect 273430 472046 273498 472102
rect 273554 472046 273622 472102
rect 273678 472046 291250 472102
rect 291306 472046 291374 472102
rect 291430 472046 291498 472102
rect 291554 472046 291622 472102
rect 291678 472046 309250 472102
rect 309306 472046 309374 472102
rect 309430 472046 309498 472102
rect 309554 472046 309622 472102
rect 309678 472046 327250 472102
rect 327306 472046 327374 472102
rect 327430 472046 327498 472102
rect 327554 472046 327622 472102
rect 327678 472046 345250 472102
rect 345306 472046 345374 472102
rect 345430 472046 345498 472102
rect 345554 472046 345622 472102
rect 345678 472046 363250 472102
rect 363306 472046 363374 472102
rect 363430 472046 363498 472102
rect 363554 472046 363622 472102
rect 363678 472046 381250 472102
rect 381306 472046 381374 472102
rect 381430 472046 381498 472102
rect 381554 472046 381622 472102
rect 381678 472046 399250 472102
rect 399306 472046 399374 472102
rect 399430 472046 399498 472102
rect 399554 472046 399622 472102
rect 399678 472046 417250 472102
rect 417306 472046 417374 472102
rect 417430 472046 417498 472102
rect 417554 472046 417622 472102
rect 417678 472046 435250 472102
rect 435306 472046 435374 472102
rect 435430 472046 435498 472102
rect 435554 472046 435622 472102
rect 435678 472046 453250 472102
rect 453306 472046 453374 472102
rect 453430 472046 453498 472102
rect 453554 472046 453622 472102
rect 453678 472046 471250 472102
rect 471306 472046 471374 472102
rect 471430 472046 471498 472102
rect 471554 472046 471622 472102
rect 471678 472046 489250 472102
rect 489306 472046 489374 472102
rect 489430 472046 489498 472102
rect 489554 472046 489622 472102
rect 489678 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 219250 471978
rect 219306 471922 219374 471978
rect 219430 471922 219498 471978
rect 219554 471922 219622 471978
rect 219678 471922 237250 471978
rect 237306 471922 237374 471978
rect 237430 471922 237498 471978
rect 237554 471922 237622 471978
rect 237678 471922 255250 471978
rect 255306 471922 255374 471978
rect 255430 471922 255498 471978
rect 255554 471922 255622 471978
rect 255678 471922 273250 471978
rect 273306 471922 273374 471978
rect 273430 471922 273498 471978
rect 273554 471922 273622 471978
rect 273678 471922 291250 471978
rect 291306 471922 291374 471978
rect 291430 471922 291498 471978
rect 291554 471922 291622 471978
rect 291678 471922 309250 471978
rect 309306 471922 309374 471978
rect 309430 471922 309498 471978
rect 309554 471922 309622 471978
rect 309678 471922 327250 471978
rect 327306 471922 327374 471978
rect 327430 471922 327498 471978
rect 327554 471922 327622 471978
rect 327678 471922 345250 471978
rect 345306 471922 345374 471978
rect 345430 471922 345498 471978
rect 345554 471922 345622 471978
rect 345678 471922 363250 471978
rect 363306 471922 363374 471978
rect 363430 471922 363498 471978
rect 363554 471922 363622 471978
rect 363678 471922 381250 471978
rect 381306 471922 381374 471978
rect 381430 471922 381498 471978
rect 381554 471922 381622 471978
rect 381678 471922 399250 471978
rect 399306 471922 399374 471978
rect 399430 471922 399498 471978
rect 399554 471922 399622 471978
rect 399678 471922 417250 471978
rect 417306 471922 417374 471978
rect 417430 471922 417498 471978
rect 417554 471922 417622 471978
rect 417678 471922 435250 471978
rect 435306 471922 435374 471978
rect 435430 471922 435498 471978
rect 435554 471922 435622 471978
rect 435678 471922 453250 471978
rect 453306 471922 453374 471978
rect 453430 471922 453498 471978
rect 453554 471922 453622 471978
rect 453678 471922 471250 471978
rect 471306 471922 471374 471978
rect 471430 471922 471498 471978
rect 471554 471922 471622 471978
rect 471678 471922 489250 471978
rect 489306 471922 489374 471978
rect 489430 471922 489498 471978
rect 489554 471922 489622 471978
rect 489678 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 204970 460350
rect 205026 460294 205094 460350
rect 205150 460294 205218 460350
rect 205274 460294 205342 460350
rect 205398 460294 222970 460350
rect 223026 460294 223094 460350
rect 223150 460294 223218 460350
rect 223274 460294 223342 460350
rect 223398 460294 240970 460350
rect 241026 460294 241094 460350
rect 241150 460294 241218 460350
rect 241274 460294 241342 460350
rect 241398 460294 258970 460350
rect 259026 460294 259094 460350
rect 259150 460294 259218 460350
rect 259274 460294 259342 460350
rect 259398 460294 276970 460350
rect 277026 460294 277094 460350
rect 277150 460294 277218 460350
rect 277274 460294 277342 460350
rect 277398 460294 294970 460350
rect 295026 460294 295094 460350
rect 295150 460294 295218 460350
rect 295274 460294 295342 460350
rect 295398 460294 312970 460350
rect 313026 460294 313094 460350
rect 313150 460294 313218 460350
rect 313274 460294 313342 460350
rect 313398 460294 330970 460350
rect 331026 460294 331094 460350
rect 331150 460294 331218 460350
rect 331274 460294 331342 460350
rect 331398 460294 348970 460350
rect 349026 460294 349094 460350
rect 349150 460294 349218 460350
rect 349274 460294 349342 460350
rect 349398 460294 366970 460350
rect 367026 460294 367094 460350
rect 367150 460294 367218 460350
rect 367274 460294 367342 460350
rect 367398 460294 384970 460350
rect 385026 460294 385094 460350
rect 385150 460294 385218 460350
rect 385274 460294 385342 460350
rect 385398 460294 402970 460350
rect 403026 460294 403094 460350
rect 403150 460294 403218 460350
rect 403274 460294 403342 460350
rect 403398 460294 420970 460350
rect 421026 460294 421094 460350
rect 421150 460294 421218 460350
rect 421274 460294 421342 460350
rect 421398 460294 438970 460350
rect 439026 460294 439094 460350
rect 439150 460294 439218 460350
rect 439274 460294 439342 460350
rect 439398 460294 456970 460350
rect 457026 460294 457094 460350
rect 457150 460294 457218 460350
rect 457274 460294 457342 460350
rect 457398 460294 474970 460350
rect 475026 460294 475094 460350
rect 475150 460294 475218 460350
rect 475274 460294 475342 460350
rect 475398 460294 492970 460350
rect 493026 460294 493094 460350
rect 493150 460294 493218 460350
rect 493274 460294 493342 460350
rect 493398 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 204970 460226
rect 205026 460170 205094 460226
rect 205150 460170 205218 460226
rect 205274 460170 205342 460226
rect 205398 460170 222970 460226
rect 223026 460170 223094 460226
rect 223150 460170 223218 460226
rect 223274 460170 223342 460226
rect 223398 460170 240970 460226
rect 241026 460170 241094 460226
rect 241150 460170 241218 460226
rect 241274 460170 241342 460226
rect 241398 460170 258970 460226
rect 259026 460170 259094 460226
rect 259150 460170 259218 460226
rect 259274 460170 259342 460226
rect 259398 460170 276970 460226
rect 277026 460170 277094 460226
rect 277150 460170 277218 460226
rect 277274 460170 277342 460226
rect 277398 460170 294970 460226
rect 295026 460170 295094 460226
rect 295150 460170 295218 460226
rect 295274 460170 295342 460226
rect 295398 460170 312970 460226
rect 313026 460170 313094 460226
rect 313150 460170 313218 460226
rect 313274 460170 313342 460226
rect 313398 460170 330970 460226
rect 331026 460170 331094 460226
rect 331150 460170 331218 460226
rect 331274 460170 331342 460226
rect 331398 460170 348970 460226
rect 349026 460170 349094 460226
rect 349150 460170 349218 460226
rect 349274 460170 349342 460226
rect 349398 460170 366970 460226
rect 367026 460170 367094 460226
rect 367150 460170 367218 460226
rect 367274 460170 367342 460226
rect 367398 460170 384970 460226
rect 385026 460170 385094 460226
rect 385150 460170 385218 460226
rect 385274 460170 385342 460226
rect 385398 460170 402970 460226
rect 403026 460170 403094 460226
rect 403150 460170 403218 460226
rect 403274 460170 403342 460226
rect 403398 460170 420970 460226
rect 421026 460170 421094 460226
rect 421150 460170 421218 460226
rect 421274 460170 421342 460226
rect 421398 460170 438970 460226
rect 439026 460170 439094 460226
rect 439150 460170 439218 460226
rect 439274 460170 439342 460226
rect 439398 460170 456970 460226
rect 457026 460170 457094 460226
rect 457150 460170 457218 460226
rect 457274 460170 457342 460226
rect 457398 460170 474970 460226
rect 475026 460170 475094 460226
rect 475150 460170 475218 460226
rect 475274 460170 475342 460226
rect 475398 460170 492970 460226
rect 493026 460170 493094 460226
rect 493150 460170 493218 460226
rect 493274 460170 493342 460226
rect 493398 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 204970 460102
rect 205026 460046 205094 460102
rect 205150 460046 205218 460102
rect 205274 460046 205342 460102
rect 205398 460046 222970 460102
rect 223026 460046 223094 460102
rect 223150 460046 223218 460102
rect 223274 460046 223342 460102
rect 223398 460046 240970 460102
rect 241026 460046 241094 460102
rect 241150 460046 241218 460102
rect 241274 460046 241342 460102
rect 241398 460046 258970 460102
rect 259026 460046 259094 460102
rect 259150 460046 259218 460102
rect 259274 460046 259342 460102
rect 259398 460046 276970 460102
rect 277026 460046 277094 460102
rect 277150 460046 277218 460102
rect 277274 460046 277342 460102
rect 277398 460046 294970 460102
rect 295026 460046 295094 460102
rect 295150 460046 295218 460102
rect 295274 460046 295342 460102
rect 295398 460046 312970 460102
rect 313026 460046 313094 460102
rect 313150 460046 313218 460102
rect 313274 460046 313342 460102
rect 313398 460046 330970 460102
rect 331026 460046 331094 460102
rect 331150 460046 331218 460102
rect 331274 460046 331342 460102
rect 331398 460046 348970 460102
rect 349026 460046 349094 460102
rect 349150 460046 349218 460102
rect 349274 460046 349342 460102
rect 349398 460046 366970 460102
rect 367026 460046 367094 460102
rect 367150 460046 367218 460102
rect 367274 460046 367342 460102
rect 367398 460046 384970 460102
rect 385026 460046 385094 460102
rect 385150 460046 385218 460102
rect 385274 460046 385342 460102
rect 385398 460046 402970 460102
rect 403026 460046 403094 460102
rect 403150 460046 403218 460102
rect 403274 460046 403342 460102
rect 403398 460046 420970 460102
rect 421026 460046 421094 460102
rect 421150 460046 421218 460102
rect 421274 460046 421342 460102
rect 421398 460046 438970 460102
rect 439026 460046 439094 460102
rect 439150 460046 439218 460102
rect 439274 460046 439342 460102
rect 439398 460046 456970 460102
rect 457026 460046 457094 460102
rect 457150 460046 457218 460102
rect 457274 460046 457342 460102
rect 457398 460046 474970 460102
rect 475026 460046 475094 460102
rect 475150 460046 475218 460102
rect 475274 460046 475342 460102
rect 475398 460046 492970 460102
rect 493026 460046 493094 460102
rect 493150 460046 493218 460102
rect 493274 460046 493342 460102
rect 493398 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 204970 459978
rect 205026 459922 205094 459978
rect 205150 459922 205218 459978
rect 205274 459922 205342 459978
rect 205398 459922 222970 459978
rect 223026 459922 223094 459978
rect 223150 459922 223218 459978
rect 223274 459922 223342 459978
rect 223398 459922 240970 459978
rect 241026 459922 241094 459978
rect 241150 459922 241218 459978
rect 241274 459922 241342 459978
rect 241398 459922 258970 459978
rect 259026 459922 259094 459978
rect 259150 459922 259218 459978
rect 259274 459922 259342 459978
rect 259398 459922 276970 459978
rect 277026 459922 277094 459978
rect 277150 459922 277218 459978
rect 277274 459922 277342 459978
rect 277398 459922 294970 459978
rect 295026 459922 295094 459978
rect 295150 459922 295218 459978
rect 295274 459922 295342 459978
rect 295398 459922 312970 459978
rect 313026 459922 313094 459978
rect 313150 459922 313218 459978
rect 313274 459922 313342 459978
rect 313398 459922 330970 459978
rect 331026 459922 331094 459978
rect 331150 459922 331218 459978
rect 331274 459922 331342 459978
rect 331398 459922 348970 459978
rect 349026 459922 349094 459978
rect 349150 459922 349218 459978
rect 349274 459922 349342 459978
rect 349398 459922 366970 459978
rect 367026 459922 367094 459978
rect 367150 459922 367218 459978
rect 367274 459922 367342 459978
rect 367398 459922 384970 459978
rect 385026 459922 385094 459978
rect 385150 459922 385218 459978
rect 385274 459922 385342 459978
rect 385398 459922 402970 459978
rect 403026 459922 403094 459978
rect 403150 459922 403218 459978
rect 403274 459922 403342 459978
rect 403398 459922 420970 459978
rect 421026 459922 421094 459978
rect 421150 459922 421218 459978
rect 421274 459922 421342 459978
rect 421398 459922 438970 459978
rect 439026 459922 439094 459978
rect 439150 459922 439218 459978
rect 439274 459922 439342 459978
rect 439398 459922 456970 459978
rect 457026 459922 457094 459978
rect 457150 459922 457218 459978
rect 457274 459922 457342 459978
rect 457398 459922 474970 459978
rect 475026 459922 475094 459978
rect 475150 459922 475218 459978
rect 475274 459922 475342 459978
rect 475398 459922 492970 459978
rect 493026 459922 493094 459978
rect 493150 459922 493218 459978
rect 493274 459922 493342 459978
rect 493398 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 165250 454350
rect 165306 454294 165374 454350
rect 165430 454294 165498 454350
rect 165554 454294 165622 454350
rect 165678 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 219250 454350
rect 219306 454294 219374 454350
rect 219430 454294 219498 454350
rect 219554 454294 219622 454350
rect 219678 454294 237250 454350
rect 237306 454294 237374 454350
rect 237430 454294 237498 454350
rect 237554 454294 237622 454350
rect 237678 454294 255250 454350
rect 255306 454294 255374 454350
rect 255430 454294 255498 454350
rect 255554 454294 255622 454350
rect 255678 454294 273250 454350
rect 273306 454294 273374 454350
rect 273430 454294 273498 454350
rect 273554 454294 273622 454350
rect 273678 454294 291250 454350
rect 291306 454294 291374 454350
rect 291430 454294 291498 454350
rect 291554 454294 291622 454350
rect 291678 454294 309250 454350
rect 309306 454294 309374 454350
rect 309430 454294 309498 454350
rect 309554 454294 309622 454350
rect 309678 454294 327250 454350
rect 327306 454294 327374 454350
rect 327430 454294 327498 454350
rect 327554 454294 327622 454350
rect 327678 454294 345250 454350
rect 345306 454294 345374 454350
rect 345430 454294 345498 454350
rect 345554 454294 345622 454350
rect 345678 454294 363250 454350
rect 363306 454294 363374 454350
rect 363430 454294 363498 454350
rect 363554 454294 363622 454350
rect 363678 454294 381250 454350
rect 381306 454294 381374 454350
rect 381430 454294 381498 454350
rect 381554 454294 381622 454350
rect 381678 454294 399250 454350
rect 399306 454294 399374 454350
rect 399430 454294 399498 454350
rect 399554 454294 399622 454350
rect 399678 454294 417250 454350
rect 417306 454294 417374 454350
rect 417430 454294 417498 454350
rect 417554 454294 417622 454350
rect 417678 454294 435250 454350
rect 435306 454294 435374 454350
rect 435430 454294 435498 454350
rect 435554 454294 435622 454350
rect 435678 454294 453250 454350
rect 453306 454294 453374 454350
rect 453430 454294 453498 454350
rect 453554 454294 453622 454350
rect 453678 454294 471250 454350
rect 471306 454294 471374 454350
rect 471430 454294 471498 454350
rect 471554 454294 471622 454350
rect 471678 454294 489250 454350
rect 489306 454294 489374 454350
rect 489430 454294 489498 454350
rect 489554 454294 489622 454350
rect 489678 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 165250 454226
rect 165306 454170 165374 454226
rect 165430 454170 165498 454226
rect 165554 454170 165622 454226
rect 165678 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 219250 454226
rect 219306 454170 219374 454226
rect 219430 454170 219498 454226
rect 219554 454170 219622 454226
rect 219678 454170 237250 454226
rect 237306 454170 237374 454226
rect 237430 454170 237498 454226
rect 237554 454170 237622 454226
rect 237678 454170 255250 454226
rect 255306 454170 255374 454226
rect 255430 454170 255498 454226
rect 255554 454170 255622 454226
rect 255678 454170 273250 454226
rect 273306 454170 273374 454226
rect 273430 454170 273498 454226
rect 273554 454170 273622 454226
rect 273678 454170 291250 454226
rect 291306 454170 291374 454226
rect 291430 454170 291498 454226
rect 291554 454170 291622 454226
rect 291678 454170 309250 454226
rect 309306 454170 309374 454226
rect 309430 454170 309498 454226
rect 309554 454170 309622 454226
rect 309678 454170 327250 454226
rect 327306 454170 327374 454226
rect 327430 454170 327498 454226
rect 327554 454170 327622 454226
rect 327678 454170 345250 454226
rect 345306 454170 345374 454226
rect 345430 454170 345498 454226
rect 345554 454170 345622 454226
rect 345678 454170 363250 454226
rect 363306 454170 363374 454226
rect 363430 454170 363498 454226
rect 363554 454170 363622 454226
rect 363678 454170 381250 454226
rect 381306 454170 381374 454226
rect 381430 454170 381498 454226
rect 381554 454170 381622 454226
rect 381678 454170 399250 454226
rect 399306 454170 399374 454226
rect 399430 454170 399498 454226
rect 399554 454170 399622 454226
rect 399678 454170 417250 454226
rect 417306 454170 417374 454226
rect 417430 454170 417498 454226
rect 417554 454170 417622 454226
rect 417678 454170 435250 454226
rect 435306 454170 435374 454226
rect 435430 454170 435498 454226
rect 435554 454170 435622 454226
rect 435678 454170 453250 454226
rect 453306 454170 453374 454226
rect 453430 454170 453498 454226
rect 453554 454170 453622 454226
rect 453678 454170 471250 454226
rect 471306 454170 471374 454226
rect 471430 454170 471498 454226
rect 471554 454170 471622 454226
rect 471678 454170 489250 454226
rect 489306 454170 489374 454226
rect 489430 454170 489498 454226
rect 489554 454170 489622 454226
rect 489678 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 165250 454102
rect 165306 454046 165374 454102
rect 165430 454046 165498 454102
rect 165554 454046 165622 454102
rect 165678 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 219250 454102
rect 219306 454046 219374 454102
rect 219430 454046 219498 454102
rect 219554 454046 219622 454102
rect 219678 454046 237250 454102
rect 237306 454046 237374 454102
rect 237430 454046 237498 454102
rect 237554 454046 237622 454102
rect 237678 454046 255250 454102
rect 255306 454046 255374 454102
rect 255430 454046 255498 454102
rect 255554 454046 255622 454102
rect 255678 454046 273250 454102
rect 273306 454046 273374 454102
rect 273430 454046 273498 454102
rect 273554 454046 273622 454102
rect 273678 454046 291250 454102
rect 291306 454046 291374 454102
rect 291430 454046 291498 454102
rect 291554 454046 291622 454102
rect 291678 454046 309250 454102
rect 309306 454046 309374 454102
rect 309430 454046 309498 454102
rect 309554 454046 309622 454102
rect 309678 454046 327250 454102
rect 327306 454046 327374 454102
rect 327430 454046 327498 454102
rect 327554 454046 327622 454102
rect 327678 454046 345250 454102
rect 345306 454046 345374 454102
rect 345430 454046 345498 454102
rect 345554 454046 345622 454102
rect 345678 454046 363250 454102
rect 363306 454046 363374 454102
rect 363430 454046 363498 454102
rect 363554 454046 363622 454102
rect 363678 454046 381250 454102
rect 381306 454046 381374 454102
rect 381430 454046 381498 454102
rect 381554 454046 381622 454102
rect 381678 454046 399250 454102
rect 399306 454046 399374 454102
rect 399430 454046 399498 454102
rect 399554 454046 399622 454102
rect 399678 454046 417250 454102
rect 417306 454046 417374 454102
rect 417430 454046 417498 454102
rect 417554 454046 417622 454102
rect 417678 454046 435250 454102
rect 435306 454046 435374 454102
rect 435430 454046 435498 454102
rect 435554 454046 435622 454102
rect 435678 454046 453250 454102
rect 453306 454046 453374 454102
rect 453430 454046 453498 454102
rect 453554 454046 453622 454102
rect 453678 454046 471250 454102
rect 471306 454046 471374 454102
rect 471430 454046 471498 454102
rect 471554 454046 471622 454102
rect 471678 454046 489250 454102
rect 489306 454046 489374 454102
rect 489430 454046 489498 454102
rect 489554 454046 489622 454102
rect 489678 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 165250 453978
rect 165306 453922 165374 453978
rect 165430 453922 165498 453978
rect 165554 453922 165622 453978
rect 165678 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 219250 453978
rect 219306 453922 219374 453978
rect 219430 453922 219498 453978
rect 219554 453922 219622 453978
rect 219678 453922 237250 453978
rect 237306 453922 237374 453978
rect 237430 453922 237498 453978
rect 237554 453922 237622 453978
rect 237678 453922 255250 453978
rect 255306 453922 255374 453978
rect 255430 453922 255498 453978
rect 255554 453922 255622 453978
rect 255678 453922 273250 453978
rect 273306 453922 273374 453978
rect 273430 453922 273498 453978
rect 273554 453922 273622 453978
rect 273678 453922 291250 453978
rect 291306 453922 291374 453978
rect 291430 453922 291498 453978
rect 291554 453922 291622 453978
rect 291678 453922 309250 453978
rect 309306 453922 309374 453978
rect 309430 453922 309498 453978
rect 309554 453922 309622 453978
rect 309678 453922 327250 453978
rect 327306 453922 327374 453978
rect 327430 453922 327498 453978
rect 327554 453922 327622 453978
rect 327678 453922 345250 453978
rect 345306 453922 345374 453978
rect 345430 453922 345498 453978
rect 345554 453922 345622 453978
rect 345678 453922 363250 453978
rect 363306 453922 363374 453978
rect 363430 453922 363498 453978
rect 363554 453922 363622 453978
rect 363678 453922 381250 453978
rect 381306 453922 381374 453978
rect 381430 453922 381498 453978
rect 381554 453922 381622 453978
rect 381678 453922 399250 453978
rect 399306 453922 399374 453978
rect 399430 453922 399498 453978
rect 399554 453922 399622 453978
rect 399678 453922 417250 453978
rect 417306 453922 417374 453978
rect 417430 453922 417498 453978
rect 417554 453922 417622 453978
rect 417678 453922 435250 453978
rect 435306 453922 435374 453978
rect 435430 453922 435498 453978
rect 435554 453922 435622 453978
rect 435678 453922 453250 453978
rect 453306 453922 453374 453978
rect 453430 453922 453498 453978
rect 453554 453922 453622 453978
rect 453678 453922 471250 453978
rect 471306 453922 471374 453978
rect 471430 453922 471498 453978
rect 471554 453922 471622 453978
rect 471678 453922 489250 453978
rect 489306 453922 489374 453978
rect 489430 453922 489498 453978
rect 489554 453922 489622 453978
rect 489678 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 114970 442350
rect 115026 442294 115094 442350
rect 115150 442294 115218 442350
rect 115274 442294 115342 442350
rect 115398 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 204970 442350
rect 205026 442294 205094 442350
rect 205150 442294 205218 442350
rect 205274 442294 205342 442350
rect 205398 442294 222970 442350
rect 223026 442294 223094 442350
rect 223150 442294 223218 442350
rect 223274 442294 223342 442350
rect 223398 442294 240970 442350
rect 241026 442294 241094 442350
rect 241150 442294 241218 442350
rect 241274 442294 241342 442350
rect 241398 442294 258970 442350
rect 259026 442294 259094 442350
rect 259150 442294 259218 442350
rect 259274 442294 259342 442350
rect 259398 442294 276970 442350
rect 277026 442294 277094 442350
rect 277150 442294 277218 442350
rect 277274 442294 277342 442350
rect 277398 442294 294970 442350
rect 295026 442294 295094 442350
rect 295150 442294 295218 442350
rect 295274 442294 295342 442350
rect 295398 442294 312970 442350
rect 313026 442294 313094 442350
rect 313150 442294 313218 442350
rect 313274 442294 313342 442350
rect 313398 442294 330970 442350
rect 331026 442294 331094 442350
rect 331150 442294 331218 442350
rect 331274 442294 331342 442350
rect 331398 442294 348970 442350
rect 349026 442294 349094 442350
rect 349150 442294 349218 442350
rect 349274 442294 349342 442350
rect 349398 442294 366970 442350
rect 367026 442294 367094 442350
rect 367150 442294 367218 442350
rect 367274 442294 367342 442350
rect 367398 442294 384970 442350
rect 385026 442294 385094 442350
rect 385150 442294 385218 442350
rect 385274 442294 385342 442350
rect 385398 442294 402970 442350
rect 403026 442294 403094 442350
rect 403150 442294 403218 442350
rect 403274 442294 403342 442350
rect 403398 442294 420970 442350
rect 421026 442294 421094 442350
rect 421150 442294 421218 442350
rect 421274 442294 421342 442350
rect 421398 442294 438970 442350
rect 439026 442294 439094 442350
rect 439150 442294 439218 442350
rect 439274 442294 439342 442350
rect 439398 442294 456970 442350
rect 457026 442294 457094 442350
rect 457150 442294 457218 442350
rect 457274 442294 457342 442350
rect 457398 442294 474970 442350
rect 475026 442294 475094 442350
rect 475150 442294 475218 442350
rect 475274 442294 475342 442350
rect 475398 442294 492970 442350
rect 493026 442294 493094 442350
rect 493150 442294 493218 442350
rect 493274 442294 493342 442350
rect 493398 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 114970 442226
rect 115026 442170 115094 442226
rect 115150 442170 115218 442226
rect 115274 442170 115342 442226
rect 115398 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 204970 442226
rect 205026 442170 205094 442226
rect 205150 442170 205218 442226
rect 205274 442170 205342 442226
rect 205398 442170 222970 442226
rect 223026 442170 223094 442226
rect 223150 442170 223218 442226
rect 223274 442170 223342 442226
rect 223398 442170 240970 442226
rect 241026 442170 241094 442226
rect 241150 442170 241218 442226
rect 241274 442170 241342 442226
rect 241398 442170 258970 442226
rect 259026 442170 259094 442226
rect 259150 442170 259218 442226
rect 259274 442170 259342 442226
rect 259398 442170 276970 442226
rect 277026 442170 277094 442226
rect 277150 442170 277218 442226
rect 277274 442170 277342 442226
rect 277398 442170 294970 442226
rect 295026 442170 295094 442226
rect 295150 442170 295218 442226
rect 295274 442170 295342 442226
rect 295398 442170 312970 442226
rect 313026 442170 313094 442226
rect 313150 442170 313218 442226
rect 313274 442170 313342 442226
rect 313398 442170 330970 442226
rect 331026 442170 331094 442226
rect 331150 442170 331218 442226
rect 331274 442170 331342 442226
rect 331398 442170 348970 442226
rect 349026 442170 349094 442226
rect 349150 442170 349218 442226
rect 349274 442170 349342 442226
rect 349398 442170 366970 442226
rect 367026 442170 367094 442226
rect 367150 442170 367218 442226
rect 367274 442170 367342 442226
rect 367398 442170 384970 442226
rect 385026 442170 385094 442226
rect 385150 442170 385218 442226
rect 385274 442170 385342 442226
rect 385398 442170 402970 442226
rect 403026 442170 403094 442226
rect 403150 442170 403218 442226
rect 403274 442170 403342 442226
rect 403398 442170 420970 442226
rect 421026 442170 421094 442226
rect 421150 442170 421218 442226
rect 421274 442170 421342 442226
rect 421398 442170 438970 442226
rect 439026 442170 439094 442226
rect 439150 442170 439218 442226
rect 439274 442170 439342 442226
rect 439398 442170 456970 442226
rect 457026 442170 457094 442226
rect 457150 442170 457218 442226
rect 457274 442170 457342 442226
rect 457398 442170 474970 442226
rect 475026 442170 475094 442226
rect 475150 442170 475218 442226
rect 475274 442170 475342 442226
rect 475398 442170 492970 442226
rect 493026 442170 493094 442226
rect 493150 442170 493218 442226
rect 493274 442170 493342 442226
rect 493398 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 114970 442102
rect 115026 442046 115094 442102
rect 115150 442046 115218 442102
rect 115274 442046 115342 442102
rect 115398 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 204970 442102
rect 205026 442046 205094 442102
rect 205150 442046 205218 442102
rect 205274 442046 205342 442102
rect 205398 442046 222970 442102
rect 223026 442046 223094 442102
rect 223150 442046 223218 442102
rect 223274 442046 223342 442102
rect 223398 442046 240970 442102
rect 241026 442046 241094 442102
rect 241150 442046 241218 442102
rect 241274 442046 241342 442102
rect 241398 442046 258970 442102
rect 259026 442046 259094 442102
rect 259150 442046 259218 442102
rect 259274 442046 259342 442102
rect 259398 442046 276970 442102
rect 277026 442046 277094 442102
rect 277150 442046 277218 442102
rect 277274 442046 277342 442102
rect 277398 442046 294970 442102
rect 295026 442046 295094 442102
rect 295150 442046 295218 442102
rect 295274 442046 295342 442102
rect 295398 442046 312970 442102
rect 313026 442046 313094 442102
rect 313150 442046 313218 442102
rect 313274 442046 313342 442102
rect 313398 442046 330970 442102
rect 331026 442046 331094 442102
rect 331150 442046 331218 442102
rect 331274 442046 331342 442102
rect 331398 442046 348970 442102
rect 349026 442046 349094 442102
rect 349150 442046 349218 442102
rect 349274 442046 349342 442102
rect 349398 442046 366970 442102
rect 367026 442046 367094 442102
rect 367150 442046 367218 442102
rect 367274 442046 367342 442102
rect 367398 442046 384970 442102
rect 385026 442046 385094 442102
rect 385150 442046 385218 442102
rect 385274 442046 385342 442102
rect 385398 442046 402970 442102
rect 403026 442046 403094 442102
rect 403150 442046 403218 442102
rect 403274 442046 403342 442102
rect 403398 442046 420970 442102
rect 421026 442046 421094 442102
rect 421150 442046 421218 442102
rect 421274 442046 421342 442102
rect 421398 442046 438970 442102
rect 439026 442046 439094 442102
rect 439150 442046 439218 442102
rect 439274 442046 439342 442102
rect 439398 442046 456970 442102
rect 457026 442046 457094 442102
rect 457150 442046 457218 442102
rect 457274 442046 457342 442102
rect 457398 442046 474970 442102
rect 475026 442046 475094 442102
rect 475150 442046 475218 442102
rect 475274 442046 475342 442102
rect 475398 442046 492970 442102
rect 493026 442046 493094 442102
rect 493150 442046 493218 442102
rect 493274 442046 493342 442102
rect 493398 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 114970 441978
rect 115026 441922 115094 441978
rect 115150 441922 115218 441978
rect 115274 441922 115342 441978
rect 115398 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 204970 441978
rect 205026 441922 205094 441978
rect 205150 441922 205218 441978
rect 205274 441922 205342 441978
rect 205398 441922 222970 441978
rect 223026 441922 223094 441978
rect 223150 441922 223218 441978
rect 223274 441922 223342 441978
rect 223398 441922 240970 441978
rect 241026 441922 241094 441978
rect 241150 441922 241218 441978
rect 241274 441922 241342 441978
rect 241398 441922 258970 441978
rect 259026 441922 259094 441978
rect 259150 441922 259218 441978
rect 259274 441922 259342 441978
rect 259398 441922 276970 441978
rect 277026 441922 277094 441978
rect 277150 441922 277218 441978
rect 277274 441922 277342 441978
rect 277398 441922 294970 441978
rect 295026 441922 295094 441978
rect 295150 441922 295218 441978
rect 295274 441922 295342 441978
rect 295398 441922 312970 441978
rect 313026 441922 313094 441978
rect 313150 441922 313218 441978
rect 313274 441922 313342 441978
rect 313398 441922 330970 441978
rect 331026 441922 331094 441978
rect 331150 441922 331218 441978
rect 331274 441922 331342 441978
rect 331398 441922 348970 441978
rect 349026 441922 349094 441978
rect 349150 441922 349218 441978
rect 349274 441922 349342 441978
rect 349398 441922 366970 441978
rect 367026 441922 367094 441978
rect 367150 441922 367218 441978
rect 367274 441922 367342 441978
rect 367398 441922 384970 441978
rect 385026 441922 385094 441978
rect 385150 441922 385218 441978
rect 385274 441922 385342 441978
rect 385398 441922 402970 441978
rect 403026 441922 403094 441978
rect 403150 441922 403218 441978
rect 403274 441922 403342 441978
rect 403398 441922 420970 441978
rect 421026 441922 421094 441978
rect 421150 441922 421218 441978
rect 421274 441922 421342 441978
rect 421398 441922 438970 441978
rect 439026 441922 439094 441978
rect 439150 441922 439218 441978
rect 439274 441922 439342 441978
rect 439398 441922 456970 441978
rect 457026 441922 457094 441978
rect 457150 441922 457218 441978
rect 457274 441922 457342 441978
rect 457398 441922 474970 441978
rect 475026 441922 475094 441978
rect 475150 441922 475218 441978
rect 475274 441922 475342 441978
rect 475398 441922 492970 441978
rect 493026 441922 493094 441978
rect 493150 441922 493218 441978
rect 493274 441922 493342 441978
rect 493398 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436378 597980 436446
rect -1916 436350 75250 436378
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436322 75250 436350
rect 75306 436322 75374 436378
rect 75430 436322 75498 436378
rect 75554 436322 75622 436378
rect 75678 436322 93250 436378
rect 93306 436322 93374 436378
rect 93430 436322 93498 436378
rect 93554 436322 93622 436378
rect 93678 436322 111250 436378
rect 111306 436322 111374 436378
rect 111430 436322 111498 436378
rect 111554 436322 111622 436378
rect 111678 436322 129250 436378
rect 129306 436322 129374 436378
rect 129430 436322 129498 436378
rect 129554 436322 129622 436378
rect 129678 436322 147250 436378
rect 147306 436322 147374 436378
rect 147430 436322 147498 436378
rect 147554 436322 147622 436378
rect 147678 436322 165250 436378
rect 165306 436322 165374 436378
rect 165430 436322 165498 436378
rect 165554 436322 165622 436378
rect 165678 436322 183250 436378
rect 183306 436322 183374 436378
rect 183430 436322 183498 436378
rect 183554 436322 183622 436378
rect 183678 436322 201250 436378
rect 201306 436322 201374 436378
rect 201430 436322 201498 436378
rect 201554 436322 201622 436378
rect 201678 436322 219250 436378
rect 219306 436322 219374 436378
rect 219430 436322 219498 436378
rect 219554 436322 219622 436378
rect 219678 436322 237250 436378
rect 237306 436322 237374 436378
rect 237430 436322 237498 436378
rect 237554 436322 237622 436378
rect 237678 436322 255250 436378
rect 255306 436322 255374 436378
rect 255430 436322 255498 436378
rect 255554 436322 255622 436378
rect 255678 436322 273250 436378
rect 273306 436322 273374 436378
rect 273430 436322 273498 436378
rect 273554 436322 273622 436378
rect 273678 436322 291250 436378
rect 291306 436322 291374 436378
rect 291430 436322 291498 436378
rect 291554 436322 291622 436378
rect 291678 436322 309250 436378
rect 309306 436322 309374 436378
rect 309430 436322 309498 436378
rect 309554 436322 309622 436378
rect 309678 436322 327250 436378
rect 327306 436322 327374 436378
rect 327430 436322 327498 436378
rect 327554 436322 327622 436378
rect 327678 436322 345250 436378
rect 345306 436322 345374 436378
rect 345430 436322 345498 436378
rect 345554 436322 345622 436378
rect 345678 436350 597980 436378
rect 345678 436322 363250 436350
rect 57678 436317 363250 436322
rect 57678 436294 64518 436317
rect -1916 436261 64518 436294
rect 64574 436261 64642 436317
rect 64698 436261 95238 436317
rect 95294 436261 95362 436317
rect 95418 436261 125958 436317
rect 126014 436261 126082 436317
rect 126138 436261 156678 436317
rect 156734 436261 156802 436317
rect 156858 436261 187398 436317
rect 187454 436261 187522 436317
rect 187578 436261 218118 436317
rect 218174 436261 218242 436317
rect 218298 436261 248838 436317
rect 248894 436261 248962 436317
rect 249018 436261 279558 436317
rect 279614 436261 279682 436317
rect 279738 436261 310278 436317
rect 310334 436261 310402 436317
rect 310458 436261 340998 436317
rect 341054 436261 341122 436317
rect 341178 436294 363250 436317
rect 363306 436294 363374 436350
rect 363430 436294 363498 436350
rect 363554 436294 363622 436350
rect 363678 436317 381250 436350
rect 363678 436294 371718 436317
rect 341178 436261 371718 436294
rect 371774 436261 371842 436317
rect 371898 436294 381250 436317
rect 381306 436294 381374 436350
rect 381430 436294 381498 436350
rect 381554 436294 381622 436350
rect 381678 436294 399250 436350
rect 399306 436294 399374 436350
rect 399430 436294 399498 436350
rect 399554 436294 399622 436350
rect 399678 436317 435250 436350
rect 399678 436294 402438 436317
rect 371898 436261 402438 436294
rect 402494 436261 402562 436317
rect 402618 436261 433158 436317
rect 433214 436261 433282 436317
rect 433338 436294 435250 436317
rect 435306 436294 435374 436350
rect 435430 436294 435498 436350
rect 435554 436294 435622 436350
rect 435678 436294 453250 436350
rect 453306 436294 453374 436350
rect 453430 436294 453498 436350
rect 453554 436294 453622 436350
rect 453678 436294 471250 436350
rect 471306 436294 471374 436350
rect 471430 436294 471498 436350
rect 471554 436294 471622 436350
rect 471678 436294 489250 436350
rect 489306 436294 489374 436350
rect 489430 436294 489498 436350
rect 489554 436294 489622 436350
rect 489678 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect 433338 436261 597980 436294
rect -1916 436254 597980 436261
rect -1916 436226 75250 436254
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436198 75250 436226
rect 75306 436198 75374 436254
rect 75430 436198 75498 436254
rect 75554 436198 75622 436254
rect 75678 436198 93250 436254
rect 93306 436198 93374 436254
rect 93430 436198 93498 436254
rect 93554 436198 93622 436254
rect 93678 436198 111250 436254
rect 111306 436198 111374 436254
rect 111430 436198 111498 436254
rect 111554 436198 111622 436254
rect 111678 436198 129250 436254
rect 129306 436198 129374 436254
rect 129430 436198 129498 436254
rect 129554 436198 129622 436254
rect 129678 436198 147250 436254
rect 147306 436198 147374 436254
rect 147430 436198 147498 436254
rect 147554 436198 147622 436254
rect 147678 436198 165250 436254
rect 165306 436198 165374 436254
rect 165430 436198 165498 436254
rect 165554 436198 165622 436254
rect 165678 436198 183250 436254
rect 183306 436198 183374 436254
rect 183430 436198 183498 436254
rect 183554 436198 183622 436254
rect 183678 436198 201250 436254
rect 201306 436198 201374 436254
rect 201430 436198 201498 436254
rect 201554 436198 201622 436254
rect 201678 436198 219250 436254
rect 219306 436198 219374 436254
rect 219430 436198 219498 436254
rect 219554 436198 219622 436254
rect 219678 436198 237250 436254
rect 237306 436198 237374 436254
rect 237430 436198 237498 436254
rect 237554 436198 237622 436254
rect 237678 436198 255250 436254
rect 255306 436198 255374 436254
rect 255430 436198 255498 436254
rect 255554 436198 255622 436254
rect 255678 436198 273250 436254
rect 273306 436198 273374 436254
rect 273430 436198 273498 436254
rect 273554 436198 273622 436254
rect 273678 436198 291250 436254
rect 291306 436198 291374 436254
rect 291430 436198 291498 436254
rect 291554 436198 291622 436254
rect 291678 436198 309250 436254
rect 309306 436198 309374 436254
rect 309430 436198 309498 436254
rect 309554 436198 309622 436254
rect 309678 436198 327250 436254
rect 327306 436198 327374 436254
rect 327430 436198 327498 436254
rect 327554 436198 327622 436254
rect 327678 436198 345250 436254
rect 345306 436198 345374 436254
rect 345430 436198 345498 436254
rect 345554 436198 345622 436254
rect 345678 436226 597980 436254
rect 345678 436198 363250 436226
rect 57678 436193 363250 436198
rect 57678 436170 64518 436193
rect -1916 436137 64518 436170
rect 64574 436137 64642 436193
rect 64698 436137 95238 436193
rect 95294 436137 95362 436193
rect 95418 436137 125958 436193
rect 126014 436137 126082 436193
rect 126138 436137 156678 436193
rect 156734 436137 156802 436193
rect 156858 436137 187398 436193
rect 187454 436137 187522 436193
rect 187578 436137 218118 436193
rect 218174 436137 218242 436193
rect 218298 436137 248838 436193
rect 248894 436137 248962 436193
rect 249018 436137 279558 436193
rect 279614 436137 279682 436193
rect 279738 436137 310278 436193
rect 310334 436137 310402 436193
rect 310458 436137 340998 436193
rect 341054 436137 341122 436193
rect 341178 436170 363250 436193
rect 363306 436170 363374 436226
rect 363430 436170 363498 436226
rect 363554 436170 363622 436226
rect 363678 436193 381250 436226
rect 363678 436170 371718 436193
rect 341178 436137 371718 436170
rect 371774 436137 371842 436193
rect 371898 436170 381250 436193
rect 381306 436170 381374 436226
rect 381430 436170 381498 436226
rect 381554 436170 381622 436226
rect 381678 436170 399250 436226
rect 399306 436170 399374 436226
rect 399430 436170 399498 436226
rect 399554 436170 399622 436226
rect 399678 436193 435250 436226
rect 399678 436170 402438 436193
rect 371898 436137 402438 436170
rect 402494 436137 402562 436193
rect 402618 436137 433158 436193
rect 433214 436137 433282 436193
rect 433338 436170 435250 436193
rect 435306 436170 435374 436226
rect 435430 436170 435498 436226
rect 435554 436170 435622 436226
rect 435678 436170 453250 436226
rect 453306 436170 453374 436226
rect 453430 436170 453498 436226
rect 453554 436170 453622 436226
rect 453678 436170 471250 436226
rect 471306 436170 471374 436226
rect 471430 436170 471498 436226
rect 471554 436170 471622 436226
rect 471678 436170 489250 436226
rect 489306 436170 489374 436226
rect 489430 436170 489498 436226
rect 489554 436170 489622 436226
rect 489678 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect 433338 436137 597980 436170
rect -1916 436130 597980 436137
rect -1916 436102 75250 436130
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436074 75250 436102
rect 75306 436074 75374 436130
rect 75430 436074 75498 436130
rect 75554 436074 75622 436130
rect 75678 436074 93250 436130
rect 93306 436074 93374 436130
rect 93430 436074 93498 436130
rect 93554 436074 93622 436130
rect 93678 436074 111250 436130
rect 111306 436074 111374 436130
rect 111430 436074 111498 436130
rect 111554 436074 111622 436130
rect 111678 436074 129250 436130
rect 129306 436074 129374 436130
rect 129430 436074 129498 436130
rect 129554 436074 129622 436130
rect 129678 436074 147250 436130
rect 147306 436074 147374 436130
rect 147430 436074 147498 436130
rect 147554 436074 147622 436130
rect 147678 436074 165250 436130
rect 165306 436074 165374 436130
rect 165430 436074 165498 436130
rect 165554 436074 165622 436130
rect 165678 436074 183250 436130
rect 183306 436074 183374 436130
rect 183430 436074 183498 436130
rect 183554 436074 183622 436130
rect 183678 436074 201250 436130
rect 201306 436074 201374 436130
rect 201430 436074 201498 436130
rect 201554 436074 201622 436130
rect 201678 436074 219250 436130
rect 219306 436074 219374 436130
rect 219430 436074 219498 436130
rect 219554 436074 219622 436130
rect 219678 436074 237250 436130
rect 237306 436074 237374 436130
rect 237430 436074 237498 436130
rect 237554 436074 237622 436130
rect 237678 436074 255250 436130
rect 255306 436074 255374 436130
rect 255430 436074 255498 436130
rect 255554 436074 255622 436130
rect 255678 436074 273250 436130
rect 273306 436074 273374 436130
rect 273430 436074 273498 436130
rect 273554 436074 273622 436130
rect 273678 436074 291250 436130
rect 291306 436074 291374 436130
rect 291430 436074 291498 436130
rect 291554 436074 291622 436130
rect 291678 436074 309250 436130
rect 309306 436074 309374 436130
rect 309430 436074 309498 436130
rect 309554 436074 309622 436130
rect 309678 436074 327250 436130
rect 327306 436074 327374 436130
rect 327430 436074 327498 436130
rect 327554 436074 327622 436130
rect 327678 436074 345250 436130
rect 345306 436074 345374 436130
rect 345430 436074 345498 436130
rect 345554 436074 345622 436130
rect 345678 436102 597980 436130
rect 345678 436074 363250 436102
rect 57678 436069 363250 436074
rect 57678 436046 64518 436069
rect -1916 436013 64518 436046
rect 64574 436013 64642 436069
rect 64698 436013 95238 436069
rect 95294 436013 95362 436069
rect 95418 436013 125958 436069
rect 126014 436013 126082 436069
rect 126138 436013 156678 436069
rect 156734 436013 156802 436069
rect 156858 436013 187398 436069
rect 187454 436013 187522 436069
rect 187578 436013 218118 436069
rect 218174 436013 218242 436069
rect 218298 436013 248838 436069
rect 248894 436013 248962 436069
rect 249018 436013 279558 436069
rect 279614 436013 279682 436069
rect 279738 436013 310278 436069
rect 310334 436013 310402 436069
rect 310458 436013 340998 436069
rect 341054 436013 341122 436069
rect 341178 436046 363250 436069
rect 363306 436046 363374 436102
rect 363430 436046 363498 436102
rect 363554 436046 363622 436102
rect 363678 436069 381250 436102
rect 363678 436046 371718 436069
rect 341178 436013 371718 436046
rect 371774 436013 371842 436069
rect 371898 436046 381250 436069
rect 381306 436046 381374 436102
rect 381430 436046 381498 436102
rect 381554 436046 381622 436102
rect 381678 436046 399250 436102
rect 399306 436046 399374 436102
rect 399430 436046 399498 436102
rect 399554 436046 399622 436102
rect 399678 436069 435250 436102
rect 399678 436046 402438 436069
rect 371898 436013 402438 436046
rect 402494 436013 402562 436069
rect 402618 436013 433158 436069
rect 433214 436013 433282 436069
rect 433338 436046 435250 436069
rect 435306 436046 435374 436102
rect 435430 436046 435498 436102
rect 435554 436046 435622 436102
rect 435678 436046 453250 436102
rect 453306 436046 453374 436102
rect 453430 436046 453498 436102
rect 453554 436046 453622 436102
rect 453678 436046 471250 436102
rect 471306 436046 471374 436102
rect 471430 436046 471498 436102
rect 471554 436046 471622 436102
rect 471678 436046 489250 436102
rect 489306 436046 489374 436102
rect 489430 436046 489498 436102
rect 489554 436046 489622 436102
rect 489678 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect 433338 436013 597980 436046
rect -1916 435978 597980 436013
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435945 363250 435978
rect 57678 435922 64518 435945
rect -1916 435889 64518 435922
rect 64574 435889 64642 435945
rect 64698 435889 95238 435945
rect 95294 435889 95362 435945
rect 95418 435889 125958 435945
rect 126014 435889 126082 435945
rect 126138 435889 156678 435945
rect 156734 435889 156802 435945
rect 156858 435889 187398 435945
rect 187454 435889 187522 435945
rect 187578 435889 218118 435945
rect 218174 435889 218242 435945
rect 218298 435889 248838 435945
rect 248894 435889 248962 435945
rect 249018 435889 279558 435945
rect 279614 435889 279682 435945
rect 279738 435889 310278 435945
rect 310334 435889 310402 435945
rect 310458 435889 340998 435945
rect 341054 435889 341122 435945
rect 341178 435922 363250 435945
rect 363306 435922 363374 435978
rect 363430 435922 363498 435978
rect 363554 435922 363622 435978
rect 363678 435945 381250 435978
rect 363678 435922 371718 435945
rect 341178 435889 371718 435922
rect 371774 435889 371842 435945
rect 371898 435922 381250 435945
rect 381306 435922 381374 435978
rect 381430 435922 381498 435978
rect 381554 435922 381622 435978
rect 381678 435922 399250 435978
rect 399306 435922 399374 435978
rect 399430 435922 399498 435978
rect 399554 435922 399622 435978
rect 399678 435945 435250 435978
rect 399678 435922 402438 435945
rect 371898 435889 402438 435922
rect 402494 435889 402562 435945
rect 402618 435889 433158 435945
rect 433214 435889 433282 435945
rect 433338 435922 435250 435945
rect 435306 435922 435374 435978
rect 435430 435922 435498 435978
rect 435554 435922 435622 435978
rect 435678 435922 453250 435978
rect 453306 435922 453374 435978
rect 453430 435922 453498 435978
rect 453554 435922 453622 435978
rect 453678 435922 471250 435978
rect 471306 435922 471374 435978
rect 471430 435922 471498 435978
rect 471554 435922 471622 435978
rect 471678 435922 489250 435978
rect 489306 435922 489374 435978
rect 489430 435922 489498 435978
rect 489554 435922 489622 435978
rect 489678 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect 433338 435889 597980 435922
rect -1916 435826 597980 435889
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 79878 424350
rect 79934 424294 80002 424350
rect 80058 424294 110598 424350
rect 110654 424294 110722 424350
rect 110778 424294 141318 424350
rect 141374 424294 141442 424350
rect 141498 424294 172038 424350
rect 172094 424294 172162 424350
rect 172218 424294 202758 424350
rect 202814 424294 202882 424350
rect 202938 424294 233478 424350
rect 233534 424294 233602 424350
rect 233658 424294 264198 424350
rect 264254 424294 264322 424350
rect 264378 424294 294918 424350
rect 294974 424294 295042 424350
rect 295098 424294 325638 424350
rect 325694 424294 325762 424350
rect 325818 424294 348970 424350
rect 349026 424294 349094 424350
rect 349150 424294 349218 424350
rect 349274 424294 349342 424350
rect 349398 424294 356358 424350
rect 356414 424294 356482 424350
rect 356538 424294 366970 424350
rect 367026 424294 367094 424350
rect 367150 424294 367218 424350
rect 367274 424294 367342 424350
rect 367398 424294 384970 424350
rect 385026 424294 385094 424350
rect 385150 424294 385218 424350
rect 385274 424294 385342 424350
rect 385398 424294 387078 424350
rect 387134 424294 387202 424350
rect 387258 424294 402970 424350
rect 403026 424294 403094 424350
rect 403150 424294 403218 424350
rect 403274 424294 403342 424350
rect 403398 424294 417798 424350
rect 417854 424294 417922 424350
rect 417978 424294 420970 424350
rect 421026 424294 421094 424350
rect 421150 424294 421218 424350
rect 421274 424294 421342 424350
rect 421398 424294 438970 424350
rect 439026 424294 439094 424350
rect 439150 424294 439218 424350
rect 439274 424294 439342 424350
rect 439398 424294 456970 424350
rect 457026 424294 457094 424350
rect 457150 424294 457218 424350
rect 457274 424294 457342 424350
rect 457398 424294 474970 424350
rect 475026 424294 475094 424350
rect 475150 424294 475218 424350
rect 475274 424294 475342 424350
rect 475398 424294 492970 424350
rect 493026 424294 493094 424350
rect 493150 424294 493218 424350
rect 493274 424294 493342 424350
rect 493398 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 79878 424226
rect 79934 424170 80002 424226
rect 80058 424170 110598 424226
rect 110654 424170 110722 424226
rect 110778 424170 141318 424226
rect 141374 424170 141442 424226
rect 141498 424170 172038 424226
rect 172094 424170 172162 424226
rect 172218 424170 202758 424226
rect 202814 424170 202882 424226
rect 202938 424170 233478 424226
rect 233534 424170 233602 424226
rect 233658 424170 264198 424226
rect 264254 424170 264322 424226
rect 264378 424170 294918 424226
rect 294974 424170 295042 424226
rect 295098 424170 325638 424226
rect 325694 424170 325762 424226
rect 325818 424170 348970 424226
rect 349026 424170 349094 424226
rect 349150 424170 349218 424226
rect 349274 424170 349342 424226
rect 349398 424170 356358 424226
rect 356414 424170 356482 424226
rect 356538 424170 366970 424226
rect 367026 424170 367094 424226
rect 367150 424170 367218 424226
rect 367274 424170 367342 424226
rect 367398 424170 384970 424226
rect 385026 424170 385094 424226
rect 385150 424170 385218 424226
rect 385274 424170 385342 424226
rect 385398 424170 387078 424226
rect 387134 424170 387202 424226
rect 387258 424170 402970 424226
rect 403026 424170 403094 424226
rect 403150 424170 403218 424226
rect 403274 424170 403342 424226
rect 403398 424170 417798 424226
rect 417854 424170 417922 424226
rect 417978 424170 420970 424226
rect 421026 424170 421094 424226
rect 421150 424170 421218 424226
rect 421274 424170 421342 424226
rect 421398 424170 438970 424226
rect 439026 424170 439094 424226
rect 439150 424170 439218 424226
rect 439274 424170 439342 424226
rect 439398 424170 456970 424226
rect 457026 424170 457094 424226
rect 457150 424170 457218 424226
rect 457274 424170 457342 424226
rect 457398 424170 474970 424226
rect 475026 424170 475094 424226
rect 475150 424170 475218 424226
rect 475274 424170 475342 424226
rect 475398 424170 492970 424226
rect 493026 424170 493094 424226
rect 493150 424170 493218 424226
rect 493274 424170 493342 424226
rect 493398 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 79878 424102
rect 79934 424046 80002 424102
rect 80058 424046 110598 424102
rect 110654 424046 110722 424102
rect 110778 424046 141318 424102
rect 141374 424046 141442 424102
rect 141498 424046 172038 424102
rect 172094 424046 172162 424102
rect 172218 424046 202758 424102
rect 202814 424046 202882 424102
rect 202938 424046 233478 424102
rect 233534 424046 233602 424102
rect 233658 424046 264198 424102
rect 264254 424046 264322 424102
rect 264378 424046 294918 424102
rect 294974 424046 295042 424102
rect 295098 424046 325638 424102
rect 325694 424046 325762 424102
rect 325818 424046 348970 424102
rect 349026 424046 349094 424102
rect 349150 424046 349218 424102
rect 349274 424046 349342 424102
rect 349398 424046 356358 424102
rect 356414 424046 356482 424102
rect 356538 424046 366970 424102
rect 367026 424046 367094 424102
rect 367150 424046 367218 424102
rect 367274 424046 367342 424102
rect 367398 424046 384970 424102
rect 385026 424046 385094 424102
rect 385150 424046 385218 424102
rect 385274 424046 385342 424102
rect 385398 424046 387078 424102
rect 387134 424046 387202 424102
rect 387258 424046 402970 424102
rect 403026 424046 403094 424102
rect 403150 424046 403218 424102
rect 403274 424046 403342 424102
rect 403398 424046 417798 424102
rect 417854 424046 417922 424102
rect 417978 424046 420970 424102
rect 421026 424046 421094 424102
rect 421150 424046 421218 424102
rect 421274 424046 421342 424102
rect 421398 424046 438970 424102
rect 439026 424046 439094 424102
rect 439150 424046 439218 424102
rect 439274 424046 439342 424102
rect 439398 424046 456970 424102
rect 457026 424046 457094 424102
rect 457150 424046 457218 424102
rect 457274 424046 457342 424102
rect 457398 424046 474970 424102
rect 475026 424046 475094 424102
rect 475150 424046 475218 424102
rect 475274 424046 475342 424102
rect 475398 424046 492970 424102
rect 493026 424046 493094 424102
rect 493150 424046 493218 424102
rect 493274 424046 493342 424102
rect 493398 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 79878 423978
rect 79934 423922 80002 423978
rect 80058 423922 110598 423978
rect 110654 423922 110722 423978
rect 110778 423922 141318 423978
rect 141374 423922 141442 423978
rect 141498 423922 172038 423978
rect 172094 423922 172162 423978
rect 172218 423922 202758 423978
rect 202814 423922 202882 423978
rect 202938 423922 233478 423978
rect 233534 423922 233602 423978
rect 233658 423922 264198 423978
rect 264254 423922 264322 423978
rect 264378 423922 294918 423978
rect 294974 423922 295042 423978
rect 295098 423922 325638 423978
rect 325694 423922 325762 423978
rect 325818 423922 348970 423978
rect 349026 423922 349094 423978
rect 349150 423922 349218 423978
rect 349274 423922 349342 423978
rect 349398 423922 356358 423978
rect 356414 423922 356482 423978
rect 356538 423922 366970 423978
rect 367026 423922 367094 423978
rect 367150 423922 367218 423978
rect 367274 423922 367342 423978
rect 367398 423922 384970 423978
rect 385026 423922 385094 423978
rect 385150 423922 385218 423978
rect 385274 423922 385342 423978
rect 385398 423922 387078 423978
rect 387134 423922 387202 423978
rect 387258 423922 402970 423978
rect 403026 423922 403094 423978
rect 403150 423922 403218 423978
rect 403274 423922 403342 423978
rect 403398 423922 417798 423978
rect 417854 423922 417922 423978
rect 417978 423922 420970 423978
rect 421026 423922 421094 423978
rect 421150 423922 421218 423978
rect 421274 423922 421342 423978
rect 421398 423922 438970 423978
rect 439026 423922 439094 423978
rect 439150 423922 439218 423978
rect 439274 423922 439342 423978
rect 439398 423922 456970 423978
rect 457026 423922 457094 423978
rect 457150 423922 457218 423978
rect 457274 423922 457342 423978
rect 457398 423922 474970 423978
rect 475026 423922 475094 423978
rect 475150 423922 475218 423978
rect 475274 423922 475342 423978
rect 475398 423922 492970 423978
rect 493026 423922 493094 423978
rect 493150 423922 493218 423978
rect 493274 423922 493342 423978
rect 493398 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 64518 418350
rect 64574 418294 64642 418350
rect 64698 418294 95238 418350
rect 95294 418294 95362 418350
rect 95418 418294 125958 418350
rect 126014 418294 126082 418350
rect 126138 418294 156678 418350
rect 156734 418294 156802 418350
rect 156858 418294 187398 418350
rect 187454 418294 187522 418350
rect 187578 418294 218118 418350
rect 218174 418294 218242 418350
rect 218298 418294 248838 418350
rect 248894 418294 248962 418350
rect 249018 418294 279558 418350
rect 279614 418294 279682 418350
rect 279738 418294 310278 418350
rect 310334 418294 310402 418350
rect 310458 418294 340998 418350
rect 341054 418294 341122 418350
rect 341178 418294 363250 418350
rect 363306 418294 363374 418350
rect 363430 418294 363498 418350
rect 363554 418294 363622 418350
rect 363678 418294 371718 418350
rect 371774 418294 371842 418350
rect 371898 418294 381250 418350
rect 381306 418294 381374 418350
rect 381430 418294 381498 418350
rect 381554 418294 381622 418350
rect 381678 418294 399250 418350
rect 399306 418294 399374 418350
rect 399430 418294 399498 418350
rect 399554 418294 399622 418350
rect 399678 418294 402438 418350
rect 402494 418294 402562 418350
rect 402618 418294 433158 418350
rect 433214 418294 433282 418350
rect 433338 418294 435250 418350
rect 435306 418294 435374 418350
rect 435430 418294 435498 418350
rect 435554 418294 435622 418350
rect 435678 418294 453250 418350
rect 453306 418294 453374 418350
rect 453430 418294 453498 418350
rect 453554 418294 453622 418350
rect 453678 418294 471250 418350
rect 471306 418294 471374 418350
rect 471430 418294 471498 418350
rect 471554 418294 471622 418350
rect 471678 418294 489250 418350
rect 489306 418294 489374 418350
rect 489430 418294 489498 418350
rect 489554 418294 489622 418350
rect 489678 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 64518 418226
rect 64574 418170 64642 418226
rect 64698 418170 95238 418226
rect 95294 418170 95362 418226
rect 95418 418170 125958 418226
rect 126014 418170 126082 418226
rect 126138 418170 156678 418226
rect 156734 418170 156802 418226
rect 156858 418170 187398 418226
rect 187454 418170 187522 418226
rect 187578 418170 218118 418226
rect 218174 418170 218242 418226
rect 218298 418170 248838 418226
rect 248894 418170 248962 418226
rect 249018 418170 279558 418226
rect 279614 418170 279682 418226
rect 279738 418170 310278 418226
rect 310334 418170 310402 418226
rect 310458 418170 340998 418226
rect 341054 418170 341122 418226
rect 341178 418170 363250 418226
rect 363306 418170 363374 418226
rect 363430 418170 363498 418226
rect 363554 418170 363622 418226
rect 363678 418170 371718 418226
rect 371774 418170 371842 418226
rect 371898 418170 381250 418226
rect 381306 418170 381374 418226
rect 381430 418170 381498 418226
rect 381554 418170 381622 418226
rect 381678 418170 399250 418226
rect 399306 418170 399374 418226
rect 399430 418170 399498 418226
rect 399554 418170 399622 418226
rect 399678 418170 402438 418226
rect 402494 418170 402562 418226
rect 402618 418170 433158 418226
rect 433214 418170 433282 418226
rect 433338 418170 435250 418226
rect 435306 418170 435374 418226
rect 435430 418170 435498 418226
rect 435554 418170 435622 418226
rect 435678 418170 453250 418226
rect 453306 418170 453374 418226
rect 453430 418170 453498 418226
rect 453554 418170 453622 418226
rect 453678 418170 471250 418226
rect 471306 418170 471374 418226
rect 471430 418170 471498 418226
rect 471554 418170 471622 418226
rect 471678 418170 489250 418226
rect 489306 418170 489374 418226
rect 489430 418170 489498 418226
rect 489554 418170 489622 418226
rect 489678 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 64518 418102
rect 64574 418046 64642 418102
rect 64698 418046 95238 418102
rect 95294 418046 95362 418102
rect 95418 418046 125958 418102
rect 126014 418046 126082 418102
rect 126138 418046 156678 418102
rect 156734 418046 156802 418102
rect 156858 418046 187398 418102
rect 187454 418046 187522 418102
rect 187578 418046 218118 418102
rect 218174 418046 218242 418102
rect 218298 418046 248838 418102
rect 248894 418046 248962 418102
rect 249018 418046 279558 418102
rect 279614 418046 279682 418102
rect 279738 418046 310278 418102
rect 310334 418046 310402 418102
rect 310458 418046 340998 418102
rect 341054 418046 341122 418102
rect 341178 418046 363250 418102
rect 363306 418046 363374 418102
rect 363430 418046 363498 418102
rect 363554 418046 363622 418102
rect 363678 418046 371718 418102
rect 371774 418046 371842 418102
rect 371898 418046 381250 418102
rect 381306 418046 381374 418102
rect 381430 418046 381498 418102
rect 381554 418046 381622 418102
rect 381678 418046 399250 418102
rect 399306 418046 399374 418102
rect 399430 418046 399498 418102
rect 399554 418046 399622 418102
rect 399678 418046 402438 418102
rect 402494 418046 402562 418102
rect 402618 418046 433158 418102
rect 433214 418046 433282 418102
rect 433338 418046 435250 418102
rect 435306 418046 435374 418102
rect 435430 418046 435498 418102
rect 435554 418046 435622 418102
rect 435678 418046 453250 418102
rect 453306 418046 453374 418102
rect 453430 418046 453498 418102
rect 453554 418046 453622 418102
rect 453678 418046 471250 418102
rect 471306 418046 471374 418102
rect 471430 418046 471498 418102
rect 471554 418046 471622 418102
rect 471678 418046 489250 418102
rect 489306 418046 489374 418102
rect 489430 418046 489498 418102
rect 489554 418046 489622 418102
rect 489678 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 64518 417978
rect 64574 417922 64642 417978
rect 64698 417922 95238 417978
rect 95294 417922 95362 417978
rect 95418 417922 125958 417978
rect 126014 417922 126082 417978
rect 126138 417922 156678 417978
rect 156734 417922 156802 417978
rect 156858 417922 187398 417978
rect 187454 417922 187522 417978
rect 187578 417922 218118 417978
rect 218174 417922 218242 417978
rect 218298 417922 248838 417978
rect 248894 417922 248962 417978
rect 249018 417922 279558 417978
rect 279614 417922 279682 417978
rect 279738 417922 310278 417978
rect 310334 417922 310402 417978
rect 310458 417922 340998 417978
rect 341054 417922 341122 417978
rect 341178 417922 363250 417978
rect 363306 417922 363374 417978
rect 363430 417922 363498 417978
rect 363554 417922 363622 417978
rect 363678 417922 371718 417978
rect 371774 417922 371842 417978
rect 371898 417922 381250 417978
rect 381306 417922 381374 417978
rect 381430 417922 381498 417978
rect 381554 417922 381622 417978
rect 381678 417922 399250 417978
rect 399306 417922 399374 417978
rect 399430 417922 399498 417978
rect 399554 417922 399622 417978
rect 399678 417922 402438 417978
rect 402494 417922 402562 417978
rect 402618 417922 433158 417978
rect 433214 417922 433282 417978
rect 433338 417922 435250 417978
rect 435306 417922 435374 417978
rect 435430 417922 435498 417978
rect 435554 417922 435622 417978
rect 435678 417922 453250 417978
rect 453306 417922 453374 417978
rect 453430 417922 453498 417978
rect 453554 417922 453622 417978
rect 453678 417922 471250 417978
rect 471306 417922 471374 417978
rect 471430 417922 471498 417978
rect 471554 417922 471622 417978
rect 471678 417922 489250 417978
rect 489306 417922 489374 417978
rect 489430 417922 489498 417978
rect 489554 417922 489622 417978
rect 489678 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 79878 406350
rect 79934 406294 80002 406350
rect 80058 406294 110598 406350
rect 110654 406294 110722 406350
rect 110778 406294 141318 406350
rect 141374 406294 141442 406350
rect 141498 406294 172038 406350
rect 172094 406294 172162 406350
rect 172218 406294 202758 406350
rect 202814 406294 202882 406350
rect 202938 406294 233478 406350
rect 233534 406294 233602 406350
rect 233658 406294 264198 406350
rect 264254 406294 264322 406350
rect 264378 406294 294918 406350
rect 294974 406294 295042 406350
rect 295098 406294 325638 406350
rect 325694 406294 325762 406350
rect 325818 406294 348970 406350
rect 349026 406294 349094 406350
rect 349150 406294 349218 406350
rect 349274 406294 349342 406350
rect 349398 406294 356358 406350
rect 356414 406294 356482 406350
rect 356538 406294 366970 406350
rect 367026 406294 367094 406350
rect 367150 406294 367218 406350
rect 367274 406294 367342 406350
rect 367398 406294 384970 406350
rect 385026 406294 385094 406350
rect 385150 406294 385218 406350
rect 385274 406294 385342 406350
rect 385398 406294 387078 406350
rect 387134 406294 387202 406350
rect 387258 406294 402970 406350
rect 403026 406294 403094 406350
rect 403150 406294 403218 406350
rect 403274 406294 403342 406350
rect 403398 406294 417798 406350
rect 417854 406294 417922 406350
rect 417978 406294 420970 406350
rect 421026 406294 421094 406350
rect 421150 406294 421218 406350
rect 421274 406294 421342 406350
rect 421398 406294 438970 406350
rect 439026 406294 439094 406350
rect 439150 406294 439218 406350
rect 439274 406294 439342 406350
rect 439398 406294 456970 406350
rect 457026 406294 457094 406350
rect 457150 406294 457218 406350
rect 457274 406294 457342 406350
rect 457398 406294 474970 406350
rect 475026 406294 475094 406350
rect 475150 406294 475218 406350
rect 475274 406294 475342 406350
rect 475398 406294 492970 406350
rect 493026 406294 493094 406350
rect 493150 406294 493218 406350
rect 493274 406294 493342 406350
rect 493398 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 79878 406226
rect 79934 406170 80002 406226
rect 80058 406170 110598 406226
rect 110654 406170 110722 406226
rect 110778 406170 141318 406226
rect 141374 406170 141442 406226
rect 141498 406170 172038 406226
rect 172094 406170 172162 406226
rect 172218 406170 202758 406226
rect 202814 406170 202882 406226
rect 202938 406170 233478 406226
rect 233534 406170 233602 406226
rect 233658 406170 264198 406226
rect 264254 406170 264322 406226
rect 264378 406170 294918 406226
rect 294974 406170 295042 406226
rect 295098 406170 325638 406226
rect 325694 406170 325762 406226
rect 325818 406170 348970 406226
rect 349026 406170 349094 406226
rect 349150 406170 349218 406226
rect 349274 406170 349342 406226
rect 349398 406170 356358 406226
rect 356414 406170 356482 406226
rect 356538 406170 366970 406226
rect 367026 406170 367094 406226
rect 367150 406170 367218 406226
rect 367274 406170 367342 406226
rect 367398 406170 384970 406226
rect 385026 406170 385094 406226
rect 385150 406170 385218 406226
rect 385274 406170 385342 406226
rect 385398 406170 387078 406226
rect 387134 406170 387202 406226
rect 387258 406170 402970 406226
rect 403026 406170 403094 406226
rect 403150 406170 403218 406226
rect 403274 406170 403342 406226
rect 403398 406170 417798 406226
rect 417854 406170 417922 406226
rect 417978 406170 420970 406226
rect 421026 406170 421094 406226
rect 421150 406170 421218 406226
rect 421274 406170 421342 406226
rect 421398 406170 438970 406226
rect 439026 406170 439094 406226
rect 439150 406170 439218 406226
rect 439274 406170 439342 406226
rect 439398 406170 456970 406226
rect 457026 406170 457094 406226
rect 457150 406170 457218 406226
rect 457274 406170 457342 406226
rect 457398 406170 474970 406226
rect 475026 406170 475094 406226
rect 475150 406170 475218 406226
rect 475274 406170 475342 406226
rect 475398 406170 492970 406226
rect 493026 406170 493094 406226
rect 493150 406170 493218 406226
rect 493274 406170 493342 406226
rect 493398 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 79878 406102
rect 79934 406046 80002 406102
rect 80058 406046 110598 406102
rect 110654 406046 110722 406102
rect 110778 406046 141318 406102
rect 141374 406046 141442 406102
rect 141498 406046 172038 406102
rect 172094 406046 172162 406102
rect 172218 406046 202758 406102
rect 202814 406046 202882 406102
rect 202938 406046 233478 406102
rect 233534 406046 233602 406102
rect 233658 406046 264198 406102
rect 264254 406046 264322 406102
rect 264378 406046 294918 406102
rect 294974 406046 295042 406102
rect 295098 406046 325638 406102
rect 325694 406046 325762 406102
rect 325818 406046 348970 406102
rect 349026 406046 349094 406102
rect 349150 406046 349218 406102
rect 349274 406046 349342 406102
rect 349398 406046 356358 406102
rect 356414 406046 356482 406102
rect 356538 406046 366970 406102
rect 367026 406046 367094 406102
rect 367150 406046 367218 406102
rect 367274 406046 367342 406102
rect 367398 406046 384970 406102
rect 385026 406046 385094 406102
rect 385150 406046 385218 406102
rect 385274 406046 385342 406102
rect 385398 406046 387078 406102
rect 387134 406046 387202 406102
rect 387258 406046 402970 406102
rect 403026 406046 403094 406102
rect 403150 406046 403218 406102
rect 403274 406046 403342 406102
rect 403398 406046 417798 406102
rect 417854 406046 417922 406102
rect 417978 406046 420970 406102
rect 421026 406046 421094 406102
rect 421150 406046 421218 406102
rect 421274 406046 421342 406102
rect 421398 406046 438970 406102
rect 439026 406046 439094 406102
rect 439150 406046 439218 406102
rect 439274 406046 439342 406102
rect 439398 406046 456970 406102
rect 457026 406046 457094 406102
rect 457150 406046 457218 406102
rect 457274 406046 457342 406102
rect 457398 406046 474970 406102
rect 475026 406046 475094 406102
rect 475150 406046 475218 406102
rect 475274 406046 475342 406102
rect 475398 406046 492970 406102
rect 493026 406046 493094 406102
rect 493150 406046 493218 406102
rect 493274 406046 493342 406102
rect 493398 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 79878 405978
rect 79934 405922 80002 405978
rect 80058 405922 110598 405978
rect 110654 405922 110722 405978
rect 110778 405922 141318 405978
rect 141374 405922 141442 405978
rect 141498 405922 172038 405978
rect 172094 405922 172162 405978
rect 172218 405922 202758 405978
rect 202814 405922 202882 405978
rect 202938 405922 233478 405978
rect 233534 405922 233602 405978
rect 233658 405922 264198 405978
rect 264254 405922 264322 405978
rect 264378 405922 294918 405978
rect 294974 405922 295042 405978
rect 295098 405922 325638 405978
rect 325694 405922 325762 405978
rect 325818 405922 348970 405978
rect 349026 405922 349094 405978
rect 349150 405922 349218 405978
rect 349274 405922 349342 405978
rect 349398 405922 356358 405978
rect 356414 405922 356482 405978
rect 356538 405922 366970 405978
rect 367026 405922 367094 405978
rect 367150 405922 367218 405978
rect 367274 405922 367342 405978
rect 367398 405922 384970 405978
rect 385026 405922 385094 405978
rect 385150 405922 385218 405978
rect 385274 405922 385342 405978
rect 385398 405922 387078 405978
rect 387134 405922 387202 405978
rect 387258 405922 402970 405978
rect 403026 405922 403094 405978
rect 403150 405922 403218 405978
rect 403274 405922 403342 405978
rect 403398 405922 417798 405978
rect 417854 405922 417922 405978
rect 417978 405922 420970 405978
rect 421026 405922 421094 405978
rect 421150 405922 421218 405978
rect 421274 405922 421342 405978
rect 421398 405922 438970 405978
rect 439026 405922 439094 405978
rect 439150 405922 439218 405978
rect 439274 405922 439342 405978
rect 439398 405922 456970 405978
rect 457026 405922 457094 405978
rect 457150 405922 457218 405978
rect 457274 405922 457342 405978
rect 457398 405922 474970 405978
rect 475026 405922 475094 405978
rect 475150 405922 475218 405978
rect 475274 405922 475342 405978
rect 475398 405922 492970 405978
rect 493026 405922 493094 405978
rect 493150 405922 493218 405978
rect 493274 405922 493342 405978
rect 493398 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 64518 400350
rect 64574 400294 64642 400350
rect 64698 400294 95238 400350
rect 95294 400294 95362 400350
rect 95418 400294 125958 400350
rect 126014 400294 126082 400350
rect 126138 400294 156678 400350
rect 156734 400294 156802 400350
rect 156858 400294 187398 400350
rect 187454 400294 187522 400350
rect 187578 400294 218118 400350
rect 218174 400294 218242 400350
rect 218298 400294 248838 400350
rect 248894 400294 248962 400350
rect 249018 400294 279558 400350
rect 279614 400294 279682 400350
rect 279738 400294 310278 400350
rect 310334 400294 310402 400350
rect 310458 400294 340998 400350
rect 341054 400294 341122 400350
rect 341178 400294 363250 400350
rect 363306 400294 363374 400350
rect 363430 400294 363498 400350
rect 363554 400294 363622 400350
rect 363678 400294 371718 400350
rect 371774 400294 371842 400350
rect 371898 400294 381250 400350
rect 381306 400294 381374 400350
rect 381430 400294 381498 400350
rect 381554 400294 381622 400350
rect 381678 400294 399250 400350
rect 399306 400294 399374 400350
rect 399430 400294 399498 400350
rect 399554 400294 399622 400350
rect 399678 400294 402438 400350
rect 402494 400294 402562 400350
rect 402618 400294 433158 400350
rect 433214 400294 433282 400350
rect 433338 400294 435250 400350
rect 435306 400294 435374 400350
rect 435430 400294 435498 400350
rect 435554 400294 435622 400350
rect 435678 400294 453250 400350
rect 453306 400294 453374 400350
rect 453430 400294 453498 400350
rect 453554 400294 453622 400350
rect 453678 400294 471250 400350
rect 471306 400294 471374 400350
rect 471430 400294 471498 400350
rect 471554 400294 471622 400350
rect 471678 400294 489250 400350
rect 489306 400294 489374 400350
rect 489430 400294 489498 400350
rect 489554 400294 489622 400350
rect 489678 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 64518 400226
rect 64574 400170 64642 400226
rect 64698 400170 95238 400226
rect 95294 400170 95362 400226
rect 95418 400170 125958 400226
rect 126014 400170 126082 400226
rect 126138 400170 156678 400226
rect 156734 400170 156802 400226
rect 156858 400170 187398 400226
rect 187454 400170 187522 400226
rect 187578 400170 218118 400226
rect 218174 400170 218242 400226
rect 218298 400170 248838 400226
rect 248894 400170 248962 400226
rect 249018 400170 279558 400226
rect 279614 400170 279682 400226
rect 279738 400170 310278 400226
rect 310334 400170 310402 400226
rect 310458 400170 340998 400226
rect 341054 400170 341122 400226
rect 341178 400170 363250 400226
rect 363306 400170 363374 400226
rect 363430 400170 363498 400226
rect 363554 400170 363622 400226
rect 363678 400170 371718 400226
rect 371774 400170 371842 400226
rect 371898 400170 381250 400226
rect 381306 400170 381374 400226
rect 381430 400170 381498 400226
rect 381554 400170 381622 400226
rect 381678 400170 399250 400226
rect 399306 400170 399374 400226
rect 399430 400170 399498 400226
rect 399554 400170 399622 400226
rect 399678 400170 402438 400226
rect 402494 400170 402562 400226
rect 402618 400170 433158 400226
rect 433214 400170 433282 400226
rect 433338 400170 435250 400226
rect 435306 400170 435374 400226
rect 435430 400170 435498 400226
rect 435554 400170 435622 400226
rect 435678 400170 453250 400226
rect 453306 400170 453374 400226
rect 453430 400170 453498 400226
rect 453554 400170 453622 400226
rect 453678 400170 471250 400226
rect 471306 400170 471374 400226
rect 471430 400170 471498 400226
rect 471554 400170 471622 400226
rect 471678 400170 489250 400226
rect 489306 400170 489374 400226
rect 489430 400170 489498 400226
rect 489554 400170 489622 400226
rect 489678 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 64518 400102
rect 64574 400046 64642 400102
rect 64698 400046 95238 400102
rect 95294 400046 95362 400102
rect 95418 400046 125958 400102
rect 126014 400046 126082 400102
rect 126138 400046 156678 400102
rect 156734 400046 156802 400102
rect 156858 400046 187398 400102
rect 187454 400046 187522 400102
rect 187578 400046 218118 400102
rect 218174 400046 218242 400102
rect 218298 400046 248838 400102
rect 248894 400046 248962 400102
rect 249018 400046 279558 400102
rect 279614 400046 279682 400102
rect 279738 400046 310278 400102
rect 310334 400046 310402 400102
rect 310458 400046 340998 400102
rect 341054 400046 341122 400102
rect 341178 400046 363250 400102
rect 363306 400046 363374 400102
rect 363430 400046 363498 400102
rect 363554 400046 363622 400102
rect 363678 400046 371718 400102
rect 371774 400046 371842 400102
rect 371898 400046 381250 400102
rect 381306 400046 381374 400102
rect 381430 400046 381498 400102
rect 381554 400046 381622 400102
rect 381678 400046 399250 400102
rect 399306 400046 399374 400102
rect 399430 400046 399498 400102
rect 399554 400046 399622 400102
rect 399678 400046 402438 400102
rect 402494 400046 402562 400102
rect 402618 400046 433158 400102
rect 433214 400046 433282 400102
rect 433338 400046 435250 400102
rect 435306 400046 435374 400102
rect 435430 400046 435498 400102
rect 435554 400046 435622 400102
rect 435678 400046 453250 400102
rect 453306 400046 453374 400102
rect 453430 400046 453498 400102
rect 453554 400046 453622 400102
rect 453678 400046 471250 400102
rect 471306 400046 471374 400102
rect 471430 400046 471498 400102
rect 471554 400046 471622 400102
rect 471678 400046 489250 400102
rect 489306 400046 489374 400102
rect 489430 400046 489498 400102
rect 489554 400046 489622 400102
rect 489678 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 64518 399978
rect 64574 399922 64642 399978
rect 64698 399922 95238 399978
rect 95294 399922 95362 399978
rect 95418 399922 125958 399978
rect 126014 399922 126082 399978
rect 126138 399922 156678 399978
rect 156734 399922 156802 399978
rect 156858 399922 187398 399978
rect 187454 399922 187522 399978
rect 187578 399922 218118 399978
rect 218174 399922 218242 399978
rect 218298 399922 248838 399978
rect 248894 399922 248962 399978
rect 249018 399922 279558 399978
rect 279614 399922 279682 399978
rect 279738 399922 310278 399978
rect 310334 399922 310402 399978
rect 310458 399922 340998 399978
rect 341054 399922 341122 399978
rect 341178 399922 363250 399978
rect 363306 399922 363374 399978
rect 363430 399922 363498 399978
rect 363554 399922 363622 399978
rect 363678 399922 371718 399978
rect 371774 399922 371842 399978
rect 371898 399922 381250 399978
rect 381306 399922 381374 399978
rect 381430 399922 381498 399978
rect 381554 399922 381622 399978
rect 381678 399922 399250 399978
rect 399306 399922 399374 399978
rect 399430 399922 399498 399978
rect 399554 399922 399622 399978
rect 399678 399922 402438 399978
rect 402494 399922 402562 399978
rect 402618 399922 433158 399978
rect 433214 399922 433282 399978
rect 433338 399922 435250 399978
rect 435306 399922 435374 399978
rect 435430 399922 435498 399978
rect 435554 399922 435622 399978
rect 435678 399922 453250 399978
rect 453306 399922 453374 399978
rect 453430 399922 453498 399978
rect 453554 399922 453622 399978
rect 453678 399922 471250 399978
rect 471306 399922 471374 399978
rect 471430 399922 471498 399978
rect 471554 399922 471622 399978
rect 471678 399922 489250 399978
rect 489306 399922 489374 399978
rect 489430 399922 489498 399978
rect 489554 399922 489622 399978
rect 489678 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 79878 388350
rect 79934 388294 80002 388350
rect 80058 388294 110598 388350
rect 110654 388294 110722 388350
rect 110778 388294 141318 388350
rect 141374 388294 141442 388350
rect 141498 388294 172038 388350
rect 172094 388294 172162 388350
rect 172218 388294 202758 388350
rect 202814 388294 202882 388350
rect 202938 388294 233478 388350
rect 233534 388294 233602 388350
rect 233658 388294 264198 388350
rect 264254 388294 264322 388350
rect 264378 388294 294918 388350
rect 294974 388294 295042 388350
rect 295098 388294 325638 388350
rect 325694 388294 325762 388350
rect 325818 388294 348970 388350
rect 349026 388294 349094 388350
rect 349150 388294 349218 388350
rect 349274 388294 349342 388350
rect 349398 388294 356358 388350
rect 356414 388294 356482 388350
rect 356538 388294 366970 388350
rect 367026 388294 367094 388350
rect 367150 388294 367218 388350
rect 367274 388294 367342 388350
rect 367398 388294 384970 388350
rect 385026 388294 385094 388350
rect 385150 388294 385218 388350
rect 385274 388294 385342 388350
rect 385398 388294 387078 388350
rect 387134 388294 387202 388350
rect 387258 388294 402970 388350
rect 403026 388294 403094 388350
rect 403150 388294 403218 388350
rect 403274 388294 403342 388350
rect 403398 388294 417798 388350
rect 417854 388294 417922 388350
rect 417978 388294 420970 388350
rect 421026 388294 421094 388350
rect 421150 388294 421218 388350
rect 421274 388294 421342 388350
rect 421398 388294 438970 388350
rect 439026 388294 439094 388350
rect 439150 388294 439218 388350
rect 439274 388294 439342 388350
rect 439398 388294 456970 388350
rect 457026 388294 457094 388350
rect 457150 388294 457218 388350
rect 457274 388294 457342 388350
rect 457398 388294 474970 388350
rect 475026 388294 475094 388350
rect 475150 388294 475218 388350
rect 475274 388294 475342 388350
rect 475398 388294 492970 388350
rect 493026 388294 493094 388350
rect 493150 388294 493218 388350
rect 493274 388294 493342 388350
rect 493398 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 79878 388226
rect 79934 388170 80002 388226
rect 80058 388170 110598 388226
rect 110654 388170 110722 388226
rect 110778 388170 141318 388226
rect 141374 388170 141442 388226
rect 141498 388170 172038 388226
rect 172094 388170 172162 388226
rect 172218 388170 202758 388226
rect 202814 388170 202882 388226
rect 202938 388170 233478 388226
rect 233534 388170 233602 388226
rect 233658 388170 264198 388226
rect 264254 388170 264322 388226
rect 264378 388170 294918 388226
rect 294974 388170 295042 388226
rect 295098 388170 325638 388226
rect 325694 388170 325762 388226
rect 325818 388170 348970 388226
rect 349026 388170 349094 388226
rect 349150 388170 349218 388226
rect 349274 388170 349342 388226
rect 349398 388170 356358 388226
rect 356414 388170 356482 388226
rect 356538 388170 366970 388226
rect 367026 388170 367094 388226
rect 367150 388170 367218 388226
rect 367274 388170 367342 388226
rect 367398 388170 384970 388226
rect 385026 388170 385094 388226
rect 385150 388170 385218 388226
rect 385274 388170 385342 388226
rect 385398 388170 387078 388226
rect 387134 388170 387202 388226
rect 387258 388170 402970 388226
rect 403026 388170 403094 388226
rect 403150 388170 403218 388226
rect 403274 388170 403342 388226
rect 403398 388170 417798 388226
rect 417854 388170 417922 388226
rect 417978 388170 420970 388226
rect 421026 388170 421094 388226
rect 421150 388170 421218 388226
rect 421274 388170 421342 388226
rect 421398 388170 438970 388226
rect 439026 388170 439094 388226
rect 439150 388170 439218 388226
rect 439274 388170 439342 388226
rect 439398 388170 456970 388226
rect 457026 388170 457094 388226
rect 457150 388170 457218 388226
rect 457274 388170 457342 388226
rect 457398 388170 474970 388226
rect 475026 388170 475094 388226
rect 475150 388170 475218 388226
rect 475274 388170 475342 388226
rect 475398 388170 492970 388226
rect 493026 388170 493094 388226
rect 493150 388170 493218 388226
rect 493274 388170 493342 388226
rect 493398 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 79878 388102
rect 79934 388046 80002 388102
rect 80058 388046 110598 388102
rect 110654 388046 110722 388102
rect 110778 388046 141318 388102
rect 141374 388046 141442 388102
rect 141498 388046 172038 388102
rect 172094 388046 172162 388102
rect 172218 388046 202758 388102
rect 202814 388046 202882 388102
rect 202938 388046 233478 388102
rect 233534 388046 233602 388102
rect 233658 388046 264198 388102
rect 264254 388046 264322 388102
rect 264378 388046 294918 388102
rect 294974 388046 295042 388102
rect 295098 388046 325638 388102
rect 325694 388046 325762 388102
rect 325818 388046 348970 388102
rect 349026 388046 349094 388102
rect 349150 388046 349218 388102
rect 349274 388046 349342 388102
rect 349398 388046 356358 388102
rect 356414 388046 356482 388102
rect 356538 388046 366970 388102
rect 367026 388046 367094 388102
rect 367150 388046 367218 388102
rect 367274 388046 367342 388102
rect 367398 388046 384970 388102
rect 385026 388046 385094 388102
rect 385150 388046 385218 388102
rect 385274 388046 385342 388102
rect 385398 388046 387078 388102
rect 387134 388046 387202 388102
rect 387258 388046 402970 388102
rect 403026 388046 403094 388102
rect 403150 388046 403218 388102
rect 403274 388046 403342 388102
rect 403398 388046 417798 388102
rect 417854 388046 417922 388102
rect 417978 388046 420970 388102
rect 421026 388046 421094 388102
rect 421150 388046 421218 388102
rect 421274 388046 421342 388102
rect 421398 388046 438970 388102
rect 439026 388046 439094 388102
rect 439150 388046 439218 388102
rect 439274 388046 439342 388102
rect 439398 388046 456970 388102
rect 457026 388046 457094 388102
rect 457150 388046 457218 388102
rect 457274 388046 457342 388102
rect 457398 388046 474970 388102
rect 475026 388046 475094 388102
rect 475150 388046 475218 388102
rect 475274 388046 475342 388102
rect 475398 388046 492970 388102
rect 493026 388046 493094 388102
rect 493150 388046 493218 388102
rect 493274 388046 493342 388102
rect 493398 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 79878 387978
rect 79934 387922 80002 387978
rect 80058 387922 110598 387978
rect 110654 387922 110722 387978
rect 110778 387922 141318 387978
rect 141374 387922 141442 387978
rect 141498 387922 172038 387978
rect 172094 387922 172162 387978
rect 172218 387922 202758 387978
rect 202814 387922 202882 387978
rect 202938 387922 233478 387978
rect 233534 387922 233602 387978
rect 233658 387922 264198 387978
rect 264254 387922 264322 387978
rect 264378 387922 294918 387978
rect 294974 387922 295042 387978
rect 295098 387922 325638 387978
rect 325694 387922 325762 387978
rect 325818 387922 348970 387978
rect 349026 387922 349094 387978
rect 349150 387922 349218 387978
rect 349274 387922 349342 387978
rect 349398 387922 356358 387978
rect 356414 387922 356482 387978
rect 356538 387922 366970 387978
rect 367026 387922 367094 387978
rect 367150 387922 367218 387978
rect 367274 387922 367342 387978
rect 367398 387922 384970 387978
rect 385026 387922 385094 387978
rect 385150 387922 385218 387978
rect 385274 387922 385342 387978
rect 385398 387922 387078 387978
rect 387134 387922 387202 387978
rect 387258 387922 402970 387978
rect 403026 387922 403094 387978
rect 403150 387922 403218 387978
rect 403274 387922 403342 387978
rect 403398 387922 417798 387978
rect 417854 387922 417922 387978
rect 417978 387922 420970 387978
rect 421026 387922 421094 387978
rect 421150 387922 421218 387978
rect 421274 387922 421342 387978
rect 421398 387922 438970 387978
rect 439026 387922 439094 387978
rect 439150 387922 439218 387978
rect 439274 387922 439342 387978
rect 439398 387922 456970 387978
rect 457026 387922 457094 387978
rect 457150 387922 457218 387978
rect 457274 387922 457342 387978
rect 457398 387922 474970 387978
rect 475026 387922 475094 387978
rect 475150 387922 475218 387978
rect 475274 387922 475342 387978
rect 475398 387922 492970 387978
rect 493026 387922 493094 387978
rect 493150 387922 493218 387978
rect 493274 387922 493342 387978
rect 493398 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 64518 382350
rect 64574 382294 64642 382350
rect 64698 382294 95238 382350
rect 95294 382294 95362 382350
rect 95418 382294 125958 382350
rect 126014 382294 126082 382350
rect 126138 382294 156678 382350
rect 156734 382294 156802 382350
rect 156858 382294 187398 382350
rect 187454 382294 187522 382350
rect 187578 382294 218118 382350
rect 218174 382294 218242 382350
rect 218298 382294 248838 382350
rect 248894 382294 248962 382350
rect 249018 382294 279558 382350
rect 279614 382294 279682 382350
rect 279738 382294 310278 382350
rect 310334 382294 310402 382350
rect 310458 382294 340998 382350
rect 341054 382294 341122 382350
rect 341178 382294 363250 382350
rect 363306 382294 363374 382350
rect 363430 382294 363498 382350
rect 363554 382294 363622 382350
rect 363678 382294 371718 382350
rect 371774 382294 371842 382350
rect 371898 382294 381250 382350
rect 381306 382294 381374 382350
rect 381430 382294 381498 382350
rect 381554 382294 381622 382350
rect 381678 382294 399250 382350
rect 399306 382294 399374 382350
rect 399430 382294 399498 382350
rect 399554 382294 399622 382350
rect 399678 382294 402438 382350
rect 402494 382294 402562 382350
rect 402618 382294 433158 382350
rect 433214 382294 433282 382350
rect 433338 382294 435250 382350
rect 435306 382294 435374 382350
rect 435430 382294 435498 382350
rect 435554 382294 435622 382350
rect 435678 382294 453250 382350
rect 453306 382294 453374 382350
rect 453430 382294 453498 382350
rect 453554 382294 453622 382350
rect 453678 382294 471250 382350
rect 471306 382294 471374 382350
rect 471430 382294 471498 382350
rect 471554 382294 471622 382350
rect 471678 382294 489250 382350
rect 489306 382294 489374 382350
rect 489430 382294 489498 382350
rect 489554 382294 489622 382350
rect 489678 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 64518 382226
rect 64574 382170 64642 382226
rect 64698 382170 95238 382226
rect 95294 382170 95362 382226
rect 95418 382170 125958 382226
rect 126014 382170 126082 382226
rect 126138 382170 156678 382226
rect 156734 382170 156802 382226
rect 156858 382170 187398 382226
rect 187454 382170 187522 382226
rect 187578 382170 218118 382226
rect 218174 382170 218242 382226
rect 218298 382170 248838 382226
rect 248894 382170 248962 382226
rect 249018 382170 279558 382226
rect 279614 382170 279682 382226
rect 279738 382170 310278 382226
rect 310334 382170 310402 382226
rect 310458 382170 340998 382226
rect 341054 382170 341122 382226
rect 341178 382170 363250 382226
rect 363306 382170 363374 382226
rect 363430 382170 363498 382226
rect 363554 382170 363622 382226
rect 363678 382170 371718 382226
rect 371774 382170 371842 382226
rect 371898 382170 381250 382226
rect 381306 382170 381374 382226
rect 381430 382170 381498 382226
rect 381554 382170 381622 382226
rect 381678 382170 399250 382226
rect 399306 382170 399374 382226
rect 399430 382170 399498 382226
rect 399554 382170 399622 382226
rect 399678 382170 402438 382226
rect 402494 382170 402562 382226
rect 402618 382170 433158 382226
rect 433214 382170 433282 382226
rect 433338 382170 435250 382226
rect 435306 382170 435374 382226
rect 435430 382170 435498 382226
rect 435554 382170 435622 382226
rect 435678 382170 453250 382226
rect 453306 382170 453374 382226
rect 453430 382170 453498 382226
rect 453554 382170 453622 382226
rect 453678 382170 471250 382226
rect 471306 382170 471374 382226
rect 471430 382170 471498 382226
rect 471554 382170 471622 382226
rect 471678 382170 489250 382226
rect 489306 382170 489374 382226
rect 489430 382170 489498 382226
rect 489554 382170 489622 382226
rect 489678 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 64518 382102
rect 64574 382046 64642 382102
rect 64698 382046 95238 382102
rect 95294 382046 95362 382102
rect 95418 382046 125958 382102
rect 126014 382046 126082 382102
rect 126138 382046 156678 382102
rect 156734 382046 156802 382102
rect 156858 382046 187398 382102
rect 187454 382046 187522 382102
rect 187578 382046 218118 382102
rect 218174 382046 218242 382102
rect 218298 382046 248838 382102
rect 248894 382046 248962 382102
rect 249018 382046 279558 382102
rect 279614 382046 279682 382102
rect 279738 382046 310278 382102
rect 310334 382046 310402 382102
rect 310458 382046 340998 382102
rect 341054 382046 341122 382102
rect 341178 382046 363250 382102
rect 363306 382046 363374 382102
rect 363430 382046 363498 382102
rect 363554 382046 363622 382102
rect 363678 382046 371718 382102
rect 371774 382046 371842 382102
rect 371898 382046 381250 382102
rect 381306 382046 381374 382102
rect 381430 382046 381498 382102
rect 381554 382046 381622 382102
rect 381678 382046 399250 382102
rect 399306 382046 399374 382102
rect 399430 382046 399498 382102
rect 399554 382046 399622 382102
rect 399678 382046 402438 382102
rect 402494 382046 402562 382102
rect 402618 382046 433158 382102
rect 433214 382046 433282 382102
rect 433338 382046 435250 382102
rect 435306 382046 435374 382102
rect 435430 382046 435498 382102
rect 435554 382046 435622 382102
rect 435678 382046 453250 382102
rect 453306 382046 453374 382102
rect 453430 382046 453498 382102
rect 453554 382046 453622 382102
rect 453678 382046 471250 382102
rect 471306 382046 471374 382102
rect 471430 382046 471498 382102
rect 471554 382046 471622 382102
rect 471678 382046 489250 382102
rect 489306 382046 489374 382102
rect 489430 382046 489498 382102
rect 489554 382046 489622 382102
rect 489678 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 64518 381978
rect 64574 381922 64642 381978
rect 64698 381922 95238 381978
rect 95294 381922 95362 381978
rect 95418 381922 125958 381978
rect 126014 381922 126082 381978
rect 126138 381922 156678 381978
rect 156734 381922 156802 381978
rect 156858 381922 187398 381978
rect 187454 381922 187522 381978
rect 187578 381922 218118 381978
rect 218174 381922 218242 381978
rect 218298 381922 248838 381978
rect 248894 381922 248962 381978
rect 249018 381922 279558 381978
rect 279614 381922 279682 381978
rect 279738 381922 310278 381978
rect 310334 381922 310402 381978
rect 310458 381922 340998 381978
rect 341054 381922 341122 381978
rect 341178 381922 363250 381978
rect 363306 381922 363374 381978
rect 363430 381922 363498 381978
rect 363554 381922 363622 381978
rect 363678 381922 371718 381978
rect 371774 381922 371842 381978
rect 371898 381922 381250 381978
rect 381306 381922 381374 381978
rect 381430 381922 381498 381978
rect 381554 381922 381622 381978
rect 381678 381922 399250 381978
rect 399306 381922 399374 381978
rect 399430 381922 399498 381978
rect 399554 381922 399622 381978
rect 399678 381922 402438 381978
rect 402494 381922 402562 381978
rect 402618 381922 433158 381978
rect 433214 381922 433282 381978
rect 433338 381922 435250 381978
rect 435306 381922 435374 381978
rect 435430 381922 435498 381978
rect 435554 381922 435622 381978
rect 435678 381922 453250 381978
rect 453306 381922 453374 381978
rect 453430 381922 453498 381978
rect 453554 381922 453622 381978
rect 453678 381922 471250 381978
rect 471306 381922 471374 381978
rect 471430 381922 471498 381978
rect 471554 381922 471622 381978
rect 471678 381922 489250 381978
rect 489306 381922 489374 381978
rect 489430 381922 489498 381978
rect 489554 381922 489622 381978
rect 489678 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 79878 370350
rect 79934 370294 80002 370350
rect 80058 370294 110598 370350
rect 110654 370294 110722 370350
rect 110778 370294 141318 370350
rect 141374 370294 141442 370350
rect 141498 370294 172038 370350
rect 172094 370294 172162 370350
rect 172218 370294 202758 370350
rect 202814 370294 202882 370350
rect 202938 370294 233478 370350
rect 233534 370294 233602 370350
rect 233658 370294 264198 370350
rect 264254 370294 264322 370350
rect 264378 370294 294918 370350
rect 294974 370294 295042 370350
rect 295098 370294 325638 370350
rect 325694 370294 325762 370350
rect 325818 370294 348970 370350
rect 349026 370294 349094 370350
rect 349150 370294 349218 370350
rect 349274 370294 349342 370350
rect 349398 370294 356358 370350
rect 356414 370294 356482 370350
rect 356538 370294 366970 370350
rect 367026 370294 367094 370350
rect 367150 370294 367218 370350
rect 367274 370294 367342 370350
rect 367398 370294 384970 370350
rect 385026 370294 385094 370350
rect 385150 370294 385218 370350
rect 385274 370294 385342 370350
rect 385398 370294 387078 370350
rect 387134 370294 387202 370350
rect 387258 370294 402970 370350
rect 403026 370294 403094 370350
rect 403150 370294 403218 370350
rect 403274 370294 403342 370350
rect 403398 370294 417798 370350
rect 417854 370294 417922 370350
rect 417978 370294 420970 370350
rect 421026 370294 421094 370350
rect 421150 370294 421218 370350
rect 421274 370294 421342 370350
rect 421398 370294 438970 370350
rect 439026 370294 439094 370350
rect 439150 370294 439218 370350
rect 439274 370294 439342 370350
rect 439398 370294 456970 370350
rect 457026 370294 457094 370350
rect 457150 370294 457218 370350
rect 457274 370294 457342 370350
rect 457398 370294 474970 370350
rect 475026 370294 475094 370350
rect 475150 370294 475218 370350
rect 475274 370294 475342 370350
rect 475398 370294 492970 370350
rect 493026 370294 493094 370350
rect 493150 370294 493218 370350
rect 493274 370294 493342 370350
rect 493398 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 79878 370226
rect 79934 370170 80002 370226
rect 80058 370170 110598 370226
rect 110654 370170 110722 370226
rect 110778 370170 141318 370226
rect 141374 370170 141442 370226
rect 141498 370170 172038 370226
rect 172094 370170 172162 370226
rect 172218 370170 202758 370226
rect 202814 370170 202882 370226
rect 202938 370170 233478 370226
rect 233534 370170 233602 370226
rect 233658 370170 264198 370226
rect 264254 370170 264322 370226
rect 264378 370170 294918 370226
rect 294974 370170 295042 370226
rect 295098 370170 325638 370226
rect 325694 370170 325762 370226
rect 325818 370170 348970 370226
rect 349026 370170 349094 370226
rect 349150 370170 349218 370226
rect 349274 370170 349342 370226
rect 349398 370170 356358 370226
rect 356414 370170 356482 370226
rect 356538 370170 366970 370226
rect 367026 370170 367094 370226
rect 367150 370170 367218 370226
rect 367274 370170 367342 370226
rect 367398 370170 384970 370226
rect 385026 370170 385094 370226
rect 385150 370170 385218 370226
rect 385274 370170 385342 370226
rect 385398 370170 387078 370226
rect 387134 370170 387202 370226
rect 387258 370170 402970 370226
rect 403026 370170 403094 370226
rect 403150 370170 403218 370226
rect 403274 370170 403342 370226
rect 403398 370170 417798 370226
rect 417854 370170 417922 370226
rect 417978 370170 420970 370226
rect 421026 370170 421094 370226
rect 421150 370170 421218 370226
rect 421274 370170 421342 370226
rect 421398 370170 438970 370226
rect 439026 370170 439094 370226
rect 439150 370170 439218 370226
rect 439274 370170 439342 370226
rect 439398 370170 456970 370226
rect 457026 370170 457094 370226
rect 457150 370170 457218 370226
rect 457274 370170 457342 370226
rect 457398 370170 474970 370226
rect 475026 370170 475094 370226
rect 475150 370170 475218 370226
rect 475274 370170 475342 370226
rect 475398 370170 492970 370226
rect 493026 370170 493094 370226
rect 493150 370170 493218 370226
rect 493274 370170 493342 370226
rect 493398 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 79878 370102
rect 79934 370046 80002 370102
rect 80058 370046 110598 370102
rect 110654 370046 110722 370102
rect 110778 370046 141318 370102
rect 141374 370046 141442 370102
rect 141498 370046 172038 370102
rect 172094 370046 172162 370102
rect 172218 370046 202758 370102
rect 202814 370046 202882 370102
rect 202938 370046 233478 370102
rect 233534 370046 233602 370102
rect 233658 370046 264198 370102
rect 264254 370046 264322 370102
rect 264378 370046 294918 370102
rect 294974 370046 295042 370102
rect 295098 370046 325638 370102
rect 325694 370046 325762 370102
rect 325818 370046 348970 370102
rect 349026 370046 349094 370102
rect 349150 370046 349218 370102
rect 349274 370046 349342 370102
rect 349398 370046 356358 370102
rect 356414 370046 356482 370102
rect 356538 370046 366970 370102
rect 367026 370046 367094 370102
rect 367150 370046 367218 370102
rect 367274 370046 367342 370102
rect 367398 370046 384970 370102
rect 385026 370046 385094 370102
rect 385150 370046 385218 370102
rect 385274 370046 385342 370102
rect 385398 370046 387078 370102
rect 387134 370046 387202 370102
rect 387258 370046 402970 370102
rect 403026 370046 403094 370102
rect 403150 370046 403218 370102
rect 403274 370046 403342 370102
rect 403398 370046 417798 370102
rect 417854 370046 417922 370102
rect 417978 370046 420970 370102
rect 421026 370046 421094 370102
rect 421150 370046 421218 370102
rect 421274 370046 421342 370102
rect 421398 370046 438970 370102
rect 439026 370046 439094 370102
rect 439150 370046 439218 370102
rect 439274 370046 439342 370102
rect 439398 370046 456970 370102
rect 457026 370046 457094 370102
rect 457150 370046 457218 370102
rect 457274 370046 457342 370102
rect 457398 370046 474970 370102
rect 475026 370046 475094 370102
rect 475150 370046 475218 370102
rect 475274 370046 475342 370102
rect 475398 370046 492970 370102
rect 493026 370046 493094 370102
rect 493150 370046 493218 370102
rect 493274 370046 493342 370102
rect 493398 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 79878 369978
rect 79934 369922 80002 369978
rect 80058 369922 110598 369978
rect 110654 369922 110722 369978
rect 110778 369922 141318 369978
rect 141374 369922 141442 369978
rect 141498 369922 172038 369978
rect 172094 369922 172162 369978
rect 172218 369922 202758 369978
rect 202814 369922 202882 369978
rect 202938 369922 233478 369978
rect 233534 369922 233602 369978
rect 233658 369922 264198 369978
rect 264254 369922 264322 369978
rect 264378 369922 294918 369978
rect 294974 369922 295042 369978
rect 295098 369922 325638 369978
rect 325694 369922 325762 369978
rect 325818 369922 348970 369978
rect 349026 369922 349094 369978
rect 349150 369922 349218 369978
rect 349274 369922 349342 369978
rect 349398 369922 356358 369978
rect 356414 369922 356482 369978
rect 356538 369922 366970 369978
rect 367026 369922 367094 369978
rect 367150 369922 367218 369978
rect 367274 369922 367342 369978
rect 367398 369922 384970 369978
rect 385026 369922 385094 369978
rect 385150 369922 385218 369978
rect 385274 369922 385342 369978
rect 385398 369922 387078 369978
rect 387134 369922 387202 369978
rect 387258 369922 402970 369978
rect 403026 369922 403094 369978
rect 403150 369922 403218 369978
rect 403274 369922 403342 369978
rect 403398 369922 417798 369978
rect 417854 369922 417922 369978
rect 417978 369922 420970 369978
rect 421026 369922 421094 369978
rect 421150 369922 421218 369978
rect 421274 369922 421342 369978
rect 421398 369922 438970 369978
rect 439026 369922 439094 369978
rect 439150 369922 439218 369978
rect 439274 369922 439342 369978
rect 439398 369922 456970 369978
rect 457026 369922 457094 369978
rect 457150 369922 457218 369978
rect 457274 369922 457342 369978
rect 457398 369922 474970 369978
rect 475026 369922 475094 369978
rect 475150 369922 475218 369978
rect 475274 369922 475342 369978
rect 475398 369922 492970 369978
rect 493026 369922 493094 369978
rect 493150 369922 493218 369978
rect 493274 369922 493342 369978
rect 493398 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 64518 364350
rect 64574 364294 64642 364350
rect 64698 364294 95238 364350
rect 95294 364294 95362 364350
rect 95418 364294 125958 364350
rect 126014 364294 126082 364350
rect 126138 364294 156678 364350
rect 156734 364294 156802 364350
rect 156858 364294 187398 364350
rect 187454 364294 187522 364350
rect 187578 364294 218118 364350
rect 218174 364294 218242 364350
rect 218298 364294 248838 364350
rect 248894 364294 248962 364350
rect 249018 364294 279558 364350
rect 279614 364294 279682 364350
rect 279738 364294 310278 364350
rect 310334 364294 310402 364350
rect 310458 364294 340998 364350
rect 341054 364294 341122 364350
rect 341178 364294 363250 364350
rect 363306 364294 363374 364350
rect 363430 364294 363498 364350
rect 363554 364294 363622 364350
rect 363678 364294 371718 364350
rect 371774 364294 371842 364350
rect 371898 364294 381250 364350
rect 381306 364294 381374 364350
rect 381430 364294 381498 364350
rect 381554 364294 381622 364350
rect 381678 364294 399250 364350
rect 399306 364294 399374 364350
rect 399430 364294 399498 364350
rect 399554 364294 399622 364350
rect 399678 364294 402438 364350
rect 402494 364294 402562 364350
rect 402618 364294 433158 364350
rect 433214 364294 433282 364350
rect 433338 364294 435250 364350
rect 435306 364294 435374 364350
rect 435430 364294 435498 364350
rect 435554 364294 435622 364350
rect 435678 364294 453250 364350
rect 453306 364294 453374 364350
rect 453430 364294 453498 364350
rect 453554 364294 453622 364350
rect 453678 364294 471250 364350
rect 471306 364294 471374 364350
rect 471430 364294 471498 364350
rect 471554 364294 471622 364350
rect 471678 364294 489250 364350
rect 489306 364294 489374 364350
rect 489430 364294 489498 364350
rect 489554 364294 489622 364350
rect 489678 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 64518 364226
rect 64574 364170 64642 364226
rect 64698 364170 95238 364226
rect 95294 364170 95362 364226
rect 95418 364170 125958 364226
rect 126014 364170 126082 364226
rect 126138 364170 156678 364226
rect 156734 364170 156802 364226
rect 156858 364170 187398 364226
rect 187454 364170 187522 364226
rect 187578 364170 218118 364226
rect 218174 364170 218242 364226
rect 218298 364170 248838 364226
rect 248894 364170 248962 364226
rect 249018 364170 279558 364226
rect 279614 364170 279682 364226
rect 279738 364170 310278 364226
rect 310334 364170 310402 364226
rect 310458 364170 340998 364226
rect 341054 364170 341122 364226
rect 341178 364170 363250 364226
rect 363306 364170 363374 364226
rect 363430 364170 363498 364226
rect 363554 364170 363622 364226
rect 363678 364170 371718 364226
rect 371774 364170 371842 364226
rect 371898 364170 381250 364226
rect 381306 364170 381374 364226
rect 381430 364170 381498 364226
rect 381554 364170 381622 364226
rect 381678 364170 399250 364226
rect 399306 364170 399374 364226
rect 399430 364170 399498 364226
rect 399554 364170 399622 364226
rect 399678 364170 402438 364226
rect 402494 364170 402562 364226
rect 402618 364170 433158 364226
rect 433214 364170 433282 364226
rect 433338 364170 435250 364226
rect 435306 364170 435374 364226
rect 435430 364170 435498 364226
rect 435554 364170 435622 364226
rect 435678 364170 453250 364226
rect 453306 364170 453374 364226
rect 453430 364170 453498 364226
rect 453554 364170 453622 364226
rect 453678 364170 471250 364226
rect 471306 364170 471374 364226
rect 471430 364170 471498 364226
rect 471554 364170 471622 364226
rect 471678 364170 489250 364226
rect 489306 364170 489374 364226
rect 489430 364170 489498 364226
rect 489554 364170 489622 364226
rect 489678 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 64518 364102
rect 64574 364046 64642 364102
rect 64698 364046 95238 364102
rect 95294 364046 95362 364102
rect 95418 364046 125958 364102
rect 126014 364046 126082 364102
rect 126138 364046 156678 364102
rect 156734 364046 156802 364102
rect 156858 364046 187398 364102
rect 187454 364046 187522 364102
rect 187578 364046 218118 364102
rect 218174 364046 218242 364102
rect 218298 364046 248838 364102
rect 248894 364046 248962 364102
rect 249018 364046 279558 364102
rect 279614 364046 279682 364102
rect 279738 364046 310278 364102
rect 310334 364046 310402 364102
rect 310458 364046 340998 364102
rect 341054 364046 341122 364102
rect 341178 364046 363250 364102
rect 363306 364046 363374 364102
rect 363430 364046 363498 364102
rect 363554 364046 363622 364102
rect 363678 364046 371718 364102
rect 371774 364046 371842 364102
rect 371898 364046 381250 364102
rect 381306 364046 381374 364102
rect 381430 364046 381498 364102
rect 381554 364046 381622 364102
rect 381678 364046 399250 364102
rect 399306 364046 399374 364102
rect 399430 364046 399498 364102
rect 399554 364046 399622 364102
rect 399678 364046 402438 364102
rect 402494 364046 402562 364102
rect 402618 364046 433158 364102
rect 433214 364046 433282 364102
rect 433338 364046 435250 364102
rect 435306 364046 435374 364102
rect 435430 364046 435498 364102
rect 435554 364046 435622 364102
rect 435678 364046 453250 364102
rect 453306 364046 453374 364102
rect 453430 364046 453498 364102
rect 453554 364046 453622 364102
rect 453678 364046 471250 364102
rect 471306 364046 471374 364102
rect 471430 364046 471498 364102
rect 471554 364046 471622 364102
rect 471678 364046 489250 364102
rect 489306 364046 489374 364102
rect 489430 364046 489498 364102
rect 489554 364046 489622 364102
rect 489678 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 64518 363978
rect 64574 363922 64642 363978
rect 64698 363922 95238 363978
rect 95294 363922 95362 363978
rect 95418 363922 125958 363978
rect 126014 363922 126082 363978
rect 126138 363922 156678 363978
rect 156734 363922 156802 363978
rect 156858 363922 187398 363978
rect 187454 363922 187522 363978
rect 187578 363922 218118 363978
rect 218174 363922 218242 363978
rect 218298 363922 248838 363978
rect 248894 363922 248962 363978
rect 249018 363922 279558 363978
rect 279614 363922 279682 363978
rect 279738 363922 310278 363978
rect 310334 363922 310402 363978
rect 310458 363922 340998 363978
rect 341054 363922 341122 363978
rect 341178 363922 363250 363978
rect 363306 363922 363374 363978
rect 363430 363922 363498 363978
rect 363554 363922 363622 363978
rect 363678 363922 371718 363978
rect 371774 363922 371842 363978
rect 371898 363922 381250 363978
rect 381306 363922 381374 363978
rect 381430 363922 381498 363978
rect 381554 363922 381622 363978
rect 381678 363922 399250 363978
rect 399306 363922 399374 363978
rect 399430 363922 399498 363978
rect 399554 363922 399622 363978
rect 399678 363922 402438 363978
rect 402494 363922 402562 363978
rect 402618 363922 433158 363978
rect 433214 363922 433282 363978
rect 433338 363922 435250 363978
rect 435306 363922 435374 363978
rect 435430 363922 435498 363978
rect 435554 363922 435622 363978
rect 435678 363922 453250 363978
rect 453306 363922 453374 363978
rect 453430 363922 453498 363978
rect 453554 363922 453622 363978
rect 453678 363922 471250 363978
rect 471306 363922 471374 363978
rect 471430 363922 471498 363978
rect 471554 363922 471622 363978
rect 471678 363922 489250 363978
rect 489306 363922 489374 363978
rect 489430 363922 489498 363978
rect 489554 363922 489622 363978
rect 489678 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 79878 352350
rect 79934 352294 80002 352350
rect 80058 352294 110598 352350
rect 110654 352294 110722 352350
rect 110778 352294 141318 352350
rect 141374 352294 141442 352350
rect 141498 352294 172038 352350
rect 172094 352294 172162 352350
rect 172218 352294 202758 352350
rect 202814 352294 202882 352350
rect 202938 352294 233478 352350
rect 233534 352294 233602 352350
rect 233658 352294 264198 352350
rect 264254 352294 264322 352350
rect 264378 352294 294918 352350
rect 294974 352294 295042 352350
rect 295098 352294 325638 352350
rect 325694 352294 325762 352350
rect 325818 352294 348970 352350
rect 349026 352294 349094 352350
rect 349150 352294 349218 352350
rect 349274 352294 349342 352350
rect 349398 352294 356358 352350
rect 356414 352294 356482 352350
rect 356538 352294 366970 352350
rect 367026 352294 367094 352350
rect 367150 352294 367218 352350
rect 367274 352294 367342 352350
rect 367398 352294 384970 352350
rect 385026 352294 385094 352350
rect 385150 352294 385218 352350
rect 385274 352294 385342 352350
rect 385398 352294 387078 352350
rect 387134 352294 387202 352350
rect 387258 352294 402970 352350
rect 403026 352294 403094 352350
rect 403150 352294 403218 352350
rect 403274 352294 403342 352350
rect 403398 352294 417798 352350
rect 417854 352294 417922 352350
rect 417978 352294 420970 352350
rect 421026 352294 421094 352350
rect 421150 352294 421218 352350
rect 421274 352294 421342 352350
rect 421398 352294 438970 352350
rect 439026 352294 439094 352350
rect 439150 352294 439218 352350
rect 439274 352294 439342 352350
rect 439398 352294 456970 352350
rect 457026 352294 457094 352350
rect 457150 352294 457218 352350
rect 457274 352294 457342 352350
rect 457398 352294 474970 352350
rect 475026 352294 475094 352350
rect 475150 352294 475218 352350
rect 475274 352294 475342 352350
rect 475398 352294 492970 352350
rect 493026 352294 493094 352350
rect 493150 352294 493218 352350
rect 493274 352294 493342 352350
rect 493398 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 79878 352226
rect 79934 352170 80002 352226
rect 80058 352170 110598 352226
rect 110654 352170 110722 352226
rect 110778 352170 141318 352226
rect 141374 352170 141442 352226
rect 141498 352170 172038 352226
rect 172094 352170 172162 352226
rect 172218 352170 202758 352226
rect 202814 352170 202882 352226
rect 202938 352170 233478 352226
rect 233534 352170 233602 352226
rect 233658 352170 264198 352226
rect 264254 352170 264322 352226
rect 264378 352170 294918 352226
rect 294974 352170 295042 352226
rect 295098 352170 325638 352226
rect 325694 352170 325762 352226
rect 325818 352170 348970 352226
rect 349026 352170 349094 352226
rect 349150 352170 349218 352226
rect 349274 352170 349342 352226
rect 349398 352170 356358 352226
rect 356414 352170 356482 352226
rect 356538 352170 366970 352226
rect 367026 352170 367094 352226
rect 367150 352170 367218 352226
rect 367274 352170 367342 352226
rect 367398 352170 384970 352226
rect 385026 352170 385094 352226
rect 385150 352170 385218 352226
rect 385274 352170 385342 352226
rect 385398 352170 387078 352226
rect 387134 352170 387202 352226
rect 387258 352170 402970 352226
rect 403026 352170 403094 352226
rect 403150 352170 403218 352226
rect 403274 352170 403342 352226
rect 403398 352170 417798 352226
rect 417854 352170 417922 352226
rect 417978 352170 420970 352226
rect 421026 352170 421094 352226
rect 421150 352170 421218 352226
rect 421274 352170 421342 352226
rect 421398 352170 438970 352226
rect 439026 352170 439094 352226
rect 439150 352170 439218 352226
rect 439274 352170 439342 352226
rect 439398 352170 456970 352226
rect 457026 352170 457094 352226
rect 457150 352170 457218 352226
rect 457274 352170 457342 352226
rect 457398 352170 474970 352226
rect 475026 352170 475094 352226
rect 475150 352170 475218 352226
rect 475274 352170 475342 352226
rect 475398 352170 492970 352226
rect 493026 352170 493094 352226
rect 493150 352170 493218 352226
rect 493274 352170 493342 352226
rect 493398 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 79878 352102
rect 79934 352046 80002 352102
rect 80058 352046 110598 352102
rect 110654 352046 110722 352102
rect 110778 352046 141318 352102
rect 141374 352046 141442 352102
rect 141498 352046 172038 352102
rect 172094 352046 172162 352102
rect 172218 352046 202758 352102
rect 202814 352046 202882 352102
rect 202938 352046 233478 352102
rect 233534 352046 233602 352102
rect 233658 352046 264198 352102
rect 264254 352046 264322 352102
rect 264378 352046 294918 352102
rect 294974 352046 295042 352102
rect 295098 352046 325638 352102
rect 325694 352046 325762 352102
rect 325818 352046 348970 352102
rect 349026 352046 349094 352102
rect 349150 352046 349218 352102
rect 349274 352046 349342 352102
rect 349398 352046 356358 352102
rect 356414 352046 356482 352102
rect 356538 352046 366970 352102
rect 367026 352046 367094 352102
rect 367150 352046 367218 352102
rect 367274 352046 367342 352102
rect 367398 352046 384970 352102
rect 385026 352046 385094 352102
rect 385150 352046 385218 352102
rect 385274 352046 385342 352102
rect 385398 352046 387078 352102
rect 387134 352046 387202 352102
rect 387258 352046 402970 352102
rect 403026 352046 403094 352102
rect 403150 352046 403218 352102
rect 403274 352046 403342 352102
rect 403398 352046 417798 352102
rect 417854 352046 417922 352102
rect 417978 352046 420970 352102
rect 421026 352046 421094 352102
rect 421150 352046 421218 352102
rect 421274 352046 421342 352102
rect 421398 352046 438970 352102
rect 439026 352046 439094 352102
rect 439150 352046 439218 352102
rect 439274 352046 439342 352102
rect 439398 352046 456970 352102
rect 457026 352046 457094 352102
rect 457150 352046 457218 352102
rect 457274 352046 457342 352102
rect 457398 352046 474970 352102
rect 475026 352046 475094 352102
rect 475150 352046 475218 352102
rect 475274 352046 475342 352102
rect 475398 352046 492970 352102
rect 493026 352046 493094 352102
rect 493150 352046 493218 352102
rect 493274 352046 493342 352102
rect 493398 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 79878 351978
rect 79934 351922 80002 351978
rect 80058 351922 110598 351978
rect 110654 351922 110722 351978
rect 110778 351922 141318 351978
rect 141374 351922 141442 351978
rect 141498 351922 172038 351978
rect 172094 351922 172162 351978
rect 172218 351922 202758 351978
rect 202814 351922 202882 351978
rect 202938 351922 233478 351978
rect 233534 351922 233602 351978
rect 233658 351922 264198 351978
rect 264254 351922 264322 351978
rect 264378 351922 294918 351978
rect 294974 351922 295042 351978
rect 295098 351922 325638 351978
rect 325694 351922 325762 351978
rect 325818 351922 348970 351978
rect 349026 351922 349094 351978
rect 349150 351922 349218 351978
rect 349274 351922 349342 351978
rect 349398 351922 356358 351978
rect 356414 351922 356482 351978
rect 356538 351922 366970 351978
rect 367026 351922 367094 351978
rect 367150 351922 367218 351978
rect 367274 351922 367342 351978
rect 367398 351922 384970 351978
rect 385026 351922 385094 351978
rect 385150 351922 385218 351978
rect 385274 351922 385342 351978
rect 385398 351922 387078 351978
rect 387134 351922 387202 351978
rect 387258 351922 402970 351978
rect 403026 351922 403094 351978
rect 403150 351922 403218 351978
rect 403274 351922 403342 351978
rect 403398 351922 417798 351978
rect 417854 351922 417922 351978
rect 417978 351922 420970 351978
rect 421026 351922 421094 351978
rect 421150 351922 421218 351978
rect 421274 351922 421342 351978
rect 421398 351922 438970 351978
rect 439026 351922 439094 351978
rect 439150 351922 439218 351978
rect 439274 351922 439342 351978
rect 439398 351922 456970 351978
rect 457026 351922 457094 351978
rect 457150 351922 457218 351978
rect 457274 351922 457342 351978
rect 457398 351922 474970 351978
rect 475026 351922 475094 351978
rect 475150 351922 475218 351978
rect 475274 351922 475342 351978
rect 475398 351922 492970 351978
rect 493026 351922 493094 351978
rect 493150 351922 493218 351978
rect 493274 351922 493342 351978
rect 493398 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 64518 346350
rect 64574 346294 64642 346350
rect 64698 346294 95238 346350
rect 95294 346294 95362 346350
rect 95418 346294 125958 346350
rect 126014 346294 126082 346350
rect 126138 346294 156678 346350
rect 156734 346294 156802 346350
rect 156858 346294 187398 346350
rect 187454 346294 187522 346350
rect 187578 346294 218118 346350
rect 218174 346294 218242 346350
rect 218298 346294 248838 346350
rect 248894 346294 248962 346350
rect 249018 346294 279558 346350
rect 279614 346294 279682 346350
rect 279738 346294 310278 346350
rect 310334 346294 310402 346350
rect 310458 346294 340998 346350
rect 341054 346294 341122 346350
rect 341178 346294 363250 346350
rect 363306 346294 363374 346350
rect 363430 346294 363498 346350
rect 363554 346294 363622 346350
rect 363678 346294 371718 346350
rect 371774 346294 371842 346350
rect 371898 346294 381250 346350
rect 381306 346294 381374 346350
rect 381430 346294 381498 346350
rect 381554 346294 381622 346350
rect 381678 346294 399250 346350
rect 399306 346294 399374 346350
rect 399430 346294 399498 346350
rect 399554 346294 399622 346350
rect 399678 346294 402438 346350
rect 402494 346294 402562 346350
rect 402618 346294 433158 346350
rect 433214 346294 433282 346350
rect 433338 346294 435250 346350
rect 435306 346294 435374 346350
rect 435430 346294 435498 346350
rect 435554 346294 435622 346350
rect 435678 346294 453250 346350
rect 453306 346294 453374 346350
rect 453430 346294 453498 346350
rect 453554 346294 453622 346350
rect 453678 346294 471250 346350
rect 471306 346294 471374 346350
rect 471430 346294 471498 346350
rect 471554 346294 471622 346350
rect 471678 346294 489250 346350
rect 489306 346294 489374 346350
rect 489430 346294 489498 346350
rect 489554 346294 489622 346350
rect 489678 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 64518 346226
rect 64574 346170 64642 346226
rect 64698 346170 95238 346226
rect 95294 346170 95362 346226
rect 95418 346170 125958 346226
rect 126014 346170 126082 346226
rect 126138 346170 156678 346226
rect 156734 346170 156802 346226
rect 156858 346170 187398 346226
rect 187454 346170 187522 346226
rect 187578 346170 218118 346226
rect 218174 346170 218242 346226
rect 218298 346170 248838 346226
rect 248894 346170 248962 346226
rect 249018 346170 279558 346226
rect 279614 346170 279682 346226
rect 279738 346170 310278 346226
rect 310334 346170 310402 346226
rect 310458 346170 340998 346226
rect 341054 346170 341122 346226
rect 341178 346170 363250 346226
rect 363306 346170 363374 346226
rect 363430 346170 363498 346226
rect 363554 346170 363622 346226
rect 363678 346170 371718 346226
rect 371774 346170 371842 346226
rect 371898 346170 381250 346226
rect 381306 346170 381374 346226
rect 381430 346170 381498 346226
rect 381554 346170 381622 346226
rect 381678 346170 399250 346226
rect 399306 346170 399374 346226
rect 399430 346170 399498 346226
rect 399554 346170 399622 346226
rect 399678 346170 402438 346226
rect 402494 346170 402562 346226
rect 402618 346170 433158 346226
rect 433214 346170 433282 346226
rect 433338 346170 435250 346226
rect 435306 346170 435374 346226
rect 435430 346170 435498 346226
rect 435554 346170 435622 346226
rect 435678 346170 453250 346226
rect 453306 346170 453374 346226
rect 453430 346170 453498 346226
rect 453554 346170 453622 346226
rect 453678 346170 471250 346226
rect 471306 346170 471374 346226
rect 471430 346170 471498 346226
rect 471554 346170 471622 346226
rect 471678 346170 489250 346226
rect 489306 346170 489374 346226
rect 489430 346170 489498 346226
rect 489554 346170 489622 346226
rect 489678 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 64518 346102
rect 64574 346046 64642 346102
rect 64698 346046 95238 346102
rect 95294 346046 95362 346102
rect 95418 346046 125958 346102
rect 126014 346046 126082 346102
rect 126138 346046 156678 346102
rect 156734 346046 156802 346102
rect 156858 346046 187398 346102
rect 187454 346046 187522 346102
rect 187578 346046 218118 346102
rect 218174 346046 218242 346102
rect 218298 346046 248838 346102
rect 248894 346046 248962 346102
rect 249018 346046 279558 346102
rect 279614 346046 279682 346102
rect 279738 346046 310278 346102
rect 310334 346046 310402 346102
rect 310458 346046 340998 346102
rect 341054 346046 341122 346102
rect 341178 346046 363250 346102
rect 363306 346046 363374 346102
rect 363430 346046 363498 346102
rect 363554 346046 363622 346102
rect 363678 346046 371718 346102
rect 371774 346046 371842 346102
rect 371898 346046 381250 346102
rect 381306 346046 381374 346102
rect 381430 346046 381498 346102
rect 381554 346046 381622 346102
rect 381678 346046 399250 346102
rect 399306 346046 399374 346102
rect 399430 346046 399498 346102
rect 399554 346046 399622 346102
rect 399678 346046 402438 346102
rect 402494 346046 402562 346102
rect 402618 346046 433158 346102
rect 433214 346046 433282 346102
rect 433338 346046 435250 346102
rect 435306 346046 435374 346102
rect 435430 346046 435498 346102
rect 435554 346046 435622 346102
rect 435678 346046 453250 346102
rect 453306 346046 453374 346102
rect 453430 346046 453498 346102
rect 453554 346046 453622 346102
rect 453678 346046 471250 346102
rect 471306 346046 471374 346102
rect 471430 346046 471498 346102
rect 471554 346046 471622 346102
rect 471678 346046 489250 346102
rect 489306 346046 489374 346102
rect 489430 346046 489498 346102
rect 489554 346046 489622 346102
rect 489678 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 64518 345978
rect 64574 345922 64642 345978
rect 64698 345922 95238 345978
rect 95294 345922 95362 345978
rect 95418 345922 125958 345978
rect 126014 345922 126082 345978
rect 126138 345922 156678 345978
rect 156734 345922 156802 345978
rect 156858 345922 187398 345978
rect 187454 345922 187522 345978
rect 187578 345922 218118 345978
rect 218174 345922 218242 345978
rect 218298 345922 248838 345978
rect 248894 345922 248962 345978
rect 249018 345922 279558 345978
rect 279614 345922 279682 345978
rect 279738 345922 310278 345978
rect 310334 345922 310402 345978
rect 310458 345922 340998 345978
rect 341054 345922 341122 345978
rect 341178 345922 363250 345978
rect 363306 345922 363374 345978
rect 363430 345922 363498 345978
rect 363554 345922 363622 345978
rect 363678 345922 371718 345978
rect 371774 345922 371842 345978
rect 371898 345922 381250 345978
rect 381306 345922 381374 345978
rect 381430 345922 381498 345978
rect 381554 345922 381622 345978
rect 381678 345922 399250 345978
rect 399306 345922 399374 345978
rect 399430 345922 399498 345978
rect 399554 345922 399622 345978
rect 399678 345922 402438 345978
rect 402494 345922 402562 345978
rect 402618 345922 433158 345978
rect 433214 345922 433282 345978
rect 433338 345922 435250 345978
rect 435306 345922 435374 345978
rect 435430 345922 435498 345978
rect 435554 345922 435622 345978
rect 435678 345922 453250 345978
rect 453306 345922 453374 345978
rect 453430 345922 453498 345978
rect 453554 345922 453622 345978
rect 453678 345922 471250 345978
rect 471306 345922 471374 345978
rect 471430 345922 471498 345978
rect 471554 345922 471622 345978
rect 471678 345922 489250 345978
rect 489306 345922 489374 345978
rect 489430 345922 489498 345978
rect 489554 345922 489622 345978
rect 489678 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 79878 334350
rect 79934 334294 80002 334350
rect 80058 334294 110598 334350
rect 110654 334294 110722 334350
rect 110778 334294 141318 334350
rect 141374 334294 141442 334350
rect 141498 334294 172038 334350
rect 172094 334294 172162 334350
rect 172218 334294 202758 334350
rect 202814 334294 202882 334350
rect 202938 334294 233478 334350
rect 233534 334294 233602 334350
rect 233658 334294 264198 334350
rect 264254 334294 264322 334350
rect 264378 334294 294918 334350
rect 294974 334294 295042 334350
rect 295098 334294 325638 334350
rect 325694 334294 325762 334350
rect 325818 334294 348970 334350
rect 349026 334294 349094 334350
rect 349150 334294 349218 334350
rect 349274 334294 349342 334350
rect 349398 334294 356358 334350
rect 356414 334294 356482 334350
rect 356538 334294 366970 334350
rect 367026 334294 367094 334350
rect 367150 334294 367218 334350
rect 367274 334294 367342 334350
rect 367398 334294 384970 334350
rect 385026 334294 385094 334350
rect 385150 334294 385218 334350
rect 385274 334294 385342 334350
rect 385398 334294 387078 334350
rect 387134 334294 387202 334350
rect 387258 334294 402970 334350
rect 403026 334294 403094 334350
rect 403150 334294 403218 334350
rect 403274 334294 403342 334350
rect 403398 334294 417798 334350
rect 417854 334294 417922 334350
rect 417978 334294 420970 334350
rect 421026 334294 421094 334350
rect 421150 334294 421218 334350
rect 421274 334294 421342 334350
rect 421398 334294 438970 334350
rect 439026 334294 439094 334350
rect 439150 334294 439218 334350
rect 439274 334294 439342 334350
rect 439398 334294 456970 334350
rect 457026 334294 457094 334350
rect 457150 334294 457218 334350
rect 457274 334294 457342 334350
rect 457398 334294 474970 334350
rect 475026 334294 475094 334350
rect 475150 334294 475218 334350
rect 475274 334294 475342 334350
rect 475398 334294 492970 334350
rect 493026 334294 493094 334350
rect 493150 334294 493218 334350
rect 493274 334294 493342 334350
rect 493398 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 79878 334226
rect 79934 334170 80002 334226
rect 80058 334170 110598 334226
rect 110654 334170 110722 334226
rect 110778 334170 141318 334226
rect 141374 334170 141442 334226
rect 141498 334170 172038 334226
rect 172094 334170 172162 334226
rect 172218 334170 202758 334226
rect 202814 334170 202882 334226
rect 202938 334170 233478 334226
rect 233534 334170 233602 334226
rect 233658 334170 264198 334226
rect 264254 334170 264322 334226
rect 264378 334170 294918 334226
rect 294974 334170 295042 334226
rect 295098 334170 325638 334226
rect 325694 334170 325762 334226
rect 325818 334170 348970 334226
rect 349026 334170 349094 334226
rect 349150 334170 349218 334226
rect 349274 334170 349342 334226
rect 349398 334170 356358 334226
rect 356414 334170 356482 334226
rect 356538 334170 366970 334226
rect 367026 334170 367094 334226
rect 367150 334170 367218 334226
rect 367274 334170 367342 334226
rect 367398 334170 384970 334226
rect 385026 334170 385094 334226
rect 385150 334170 385218 334226
rect 385274 334170 385342 334226
rect 385398 334170 387078 334226
rect 387134 334170 387202 334226
rect 387258 334170 402970 334226
rect 403026 334170 403094 334226
rect 403150 334170 403218 334226
rect 403274 334170 403342 334226
rect 403398 334170 417798 334226
rect 417854 334170 417922 334226
rect 417978 334170 420970 334226
rect 421026 334170 421094 334226
rect 421150 334170 421218 334226
rect 421274 334170 421342 334226
rect 421398 334170 438970 334226
rect 439026 334170 439094 334226
rect 439150 334170 439218 334226
rect 439274 334170 439342 334226
rect 439398 334170 456970 334226
rect 457026 334170 457094 334226
rect 457150 334170 457218 334226
rect 457274 334170 457342 334226
rect 457398 334170 474970 334226
rect 475026 334170 475094 334226
rect 475150 334170 475218 334226
rect 475274 334170 475342 334226
rect 475398 334170 492970 334226
rect 493026 334170 493094 334226
rect 493150 334170 493218 334226
rect 493274 334170 493342 334226
rect 493398 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 79878 334102
rect 79934 334046 80002 334102
rect 80058 334046 110598 334102
rect 110654 334046 110722 334102
rect 110778 334046 141318 334102
rect 141374 334046 141442 334102
rect 141498 334046 172038 334102
rect 172094 334046 172162 334102
rect 172218 334046 202758 334102
rect 202814 334046 202882 334102
rect 202938 334046 233478 334102
rect 233534 334046 233602 334102
rect 233658 334046 264198 334102
rect 264254 334046 264322 334102
rect 264378 334046 294918 334102
rect 294974 334046 295042 334102
rect 295098 334046 325638 334102
rect 325694 334046 325762 334102
rect 325818 334046 348970 334102
rect 349026 334046 349094 334102
rect 349150 334046 349218 334102
rect 349274 334046 349342 334102
rect 349398 334046 356358 334102
rect 356414 334046 356482 334102
rect 356538 334046 366970 334102
rect 367026 334046 367094 334102
rect 367150 334046 367218 334102
rect 367274 334046 367342 334102
rect 367398 334046 384970 334102
rect 385026 334046 385094 334102
rect 385150 334046 385218 334102
rect 385274 334046 385342 334102
rect 385398 334046 387078 334102
rect 387134 334046 387202 334102
rect 387258 334046 402970 334102
rect 403026 334046 403094 334102
rect 403150 334046 403218 334102
rect 403274 334046 403342 334102
rect 403398 334046 417798 334102
rect 417854 334046 417922 334102
rect 417978 334046 420970 334102
rect 421026 334046 421094 334102
rect 421150 334046 421218 334102
rect 421274 334046 421342 334102
rect 421398 334046 438970 334102
rect 439026 334046 439094 334102
rect 439150 334046 439218 334102
rect 439274 334046 439342 334102
rect 439398 334046 456970 334102
rect 457026 334046 457094 334102
rect 457150 334046 457218 334102
rect 457274 334046 457342 334102
rect 457398 334046 474970 334102
rect 475026 334046 475094 334102
rect 475150 334046 475218 334102
rect 475274 334046 475342 334102
rect 475398 334046 492970 334102
rect 493026 334046 493094 334102
rect 493150 334046 493218 334102
rect 493274 334046 493342 334102
rect 493398 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 79878 333978
rect 79934 333922 80002 333978
rect 80058 333922 110598 333978
rect 110654 333922 110722 333978
rect 110778 333922 141318 333978
rect 141374 333922 141442 333978
rect 141498 333922 172038 333978
rect 172094 333922 172162 333978
rect 172218 333922 202758 333978
rect 202814 333922 202882 333978
rect 202938 333922 233478 333978
rect 233534 333922 233602 333978
rect 233658 333922 264198 333978
rect 264254 333922 264322 333978
rect 264378 333922 294918 333978
rect 294974 333922 295042 333978
rect 295098 333922 325638 333978
rect 325694 333922 325762 333978
rect 325818 333922 348970 333978
rect 349026 333922 349094 333978
rect 349150 333922 349218 333978
rect 349274 333922 349342 333978
rect 349398 333922 356358 333978
rect 356414 333922 356482 333978
rect 356538 333922 366970 333978
rect 367026 333922 367094 333978
rect 367150 333922 367218 333978
rect 367274 333922 367342 333978
rect 367398 333922 384970 333978
rect 385026 333922 385094 333978
rect 385150 333922 385218 333978
rect 385274 333922 385342 333978
rect 385398 333922 387078 333978
rect 387134 333922 387202 333978
rect 387258 333922 402970 333978
rect 403026 333922 403094 333978
rect 403150 333922 403218 333978
rect 403274 333922 403342 333978
rect 403398 333922 417798 333978
rect 417854 333922 417922 333978
rect 417978 333922 420970 333978
rect 421026 333922 421094 333978
rect 421150 333922 421218 333978
rect 421274 333922 421342 333978
rect 421398 333922 438970 333978
rect 439026 333922 439094 333978
rect 439150 333922 439218 333978
rect 439274 333922 439342 333978
rect 439398 333922 456970 333978
rect 457026 333922 457094 333978
rect 457150 333922 457218 333978
rect 457274 333922 457342 333978
rect 457398 333922 474970 333978
rect 475026 333922 475094 333978
rect 475150 333922 475218 333978
rect 475274 333922 475342 333978
rect 475398 333922 492970 333978
rect 493026 333922 493094 333978
rect 493150 333922 493218 333978
rect 493274 333922 493342 333978
rect 493398 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 64518 328350
rect 64574 328294 64642 328350
rect 64698 328294 95238 328350
rect 95294 328294 95362 328350
rect 95418 328294 125958 328350
rect 126014 328294 126082 328350
rect 126138 328294 156678 328350
rect 156734 328294 156802 328350
rect 156858 328294 187398 328350
rect 187454 328294 187522 328350
rect 187578 328294 218118 328350
rect 218174 328294 218242 328350
rect 218298 328294 248838 328350
rect 248894 328294 248962 328350
rect 249018 328294 279558 328350
rect 279614 328294 279682 328350
rect 279738 328294 310278 328350
rect 310334 328294 310402 328350
rect 310458 328294 340998 328350
rect 341054 328294 341122 328350
rect 341178 328294 363250 328350
rect 363306 328294 363374 328350
rect 363430 328294 363498 328350
rect 363554 328294 363622 328350
rect 363678 328294 371718 328350
rect 371774 328294 371842 328350
rect 371898 328294 381250 328350
rect 381306 328294 381374 328350
rect 381430 328294 381498 328350
rect 381554 328294 381622 328350
rect 381678 328294 399250 328350
rect 399306 328294 399374 328350
rect 399430 328294 399498 328350
rect 399554 328294 399622 328350
rect 399678 328294 402438 328350
rect 402494 328294 402562 328350
rect 402618 328294 433158 328350
rect 433214 328294 433282 328350
rect 433338 328294 435250 328350
rect 435306 328294 435374 328350
rect 435430 328294 435498 328350
rect 435554 328294 435622 328350
rect 435678 328294 453250 328350
rect 453306 328294 453374 328350
rect 453430 328294 453498 328350
rect 453554 328294 453622 328350
rect 453678 328294 471250 328350
rect 471306 328294 471374 328350
rect 471430 328294 471498 328350
rect 471554 328294 471622 328350
rect 471678 328294 489250 328350
rect 489306 328294 489374 328350
rect 489430 328294 489498 328350
rect 489554 328294 489622 328350
rect 489678 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 64518 328226
rect 64574 328170 64642 328226
rect 64698 328170 95238 328226
rect 95294 328170 95362 328226
rect 95418 328170 125958 328226
rect 126014 328170 126082 328226
rect 126138 328170 156678 328226
rect 156734 328170 156802 328226
rect 156858 328170 187398 328226
rect 187454 328170 187522 328226
rect 187578 328170 218118 328226
rect 218174 328170 218242 328226
rect 218298 328170 248838 328226
rect 248894 328170 248962 328226
rect 249018 328170 279558 328226
rect 279614 328170 279682 328226
rect 279738 328170 310278 328226
rect 310334 328170 310402 328226
rect 310458 328170 340998 328226
rect 341054 328170 341122 328226
rect 341178 328170 363250 328226
rect 363306 328170 363374 328226
rect 363430 328170 363498 328226
rect 363554 328170 363622 328226
rect 363678 328170 371718 328226
rect 371774 328170 371842 328226
rect 371898 328170 381250 328226
rect 381306 328170 381374 328226
rect 381430 328170 381498 328226
rect 381554 328170 381622 328226
rect 381678 328170 399250 328226
rect 399306 328170 399374 328226
rect 399430 328170 399498 328226
rect 399554 328170 399622 328226
rect 399678 328170 402438 328226
rect 402494 328170 402562 328226
rect 402618 328170 433158 328226
rect 433214 328170 433282 328226
rect 433338 328170 435250 328226
rect 435306 328170 435374 328226
rect 435430 328170 435498 328226
rect 435554 328170 435622 328226
rect 435678 328170 453250 328226
rect 453306 328170 453374 328226
rect 453430 328170 453498 328226
rect 453554 328170 453622 328226
rect 453678 328170 471250 328226
rect 471306 328170 471374 328226
rect 471430 328170 471498 328226
rect 471554 328170 471622 328226
rect 471678 328170 489250 328226
rect 489306 328170 489374 328226
rect 489430 328170 489498 328226
rect 489554 328170 489622 328226
rect 489678 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 64518 328102
rect 64574 328046 64642 328102
rect 64698 328046 95238 328102
rect 95294 328046 95362 328102
rect 95418 328046 125958 328102
rect 126014 328046 126082 328102
rect 126138 328046 156678 328102
rect 156734 328046 156802 328102
rect 156858 328046 187398 328102
rect 187454 328046 187522 328102
rect 187578 328046 218118 328102
rect 218174 328046 218242 328102
rect 218298 328046 248838 328102
rect 248894 328046 248962 328102
rect 249018 328046 279558 328102
rect 279614 328046 279682 328102
rect 279738 328046 310278 328102
rect 310334 328046 310402 328102
rect 310458 328046 340998 328102
rect 341054 328046 341122 328102
rect 341178 328046 363250 328102
rect 363306 328046 363374 328102
rect 363430 328046 363498 328102
rect 363554 328046 363622 328102
rect 363678 328046 371718 328102
rect 371774 328046 371842 328102
rect 371898 328046 381250 328102
rect 381306 328046 381374 328102
rect 381430 328046 381498 328102
rect 381554 328046 381622 328102
rect 381678 328046 399250 328102
rect 399306 328046 399374 328102
rect 399430 328046 399498 328102
rect 399554 328046 399622 328102
rect 399678 328046 402438 328102
rect 402494 328046 402562 328102
rect 402618 328046 433158 328102
rect 433214 328046 433282 328102
rect 433338 328046 435250 328102
rect 435306 328046 435374 328102
rect 435430 328046 435498 328102
rect 435554 328046 435622 328102
rect 435678 328046 453250 328102
rect 453306 328046 453374 328102
rect 453430 328046 453498 328102
rect 453554 328046 453622 328102
rect 453678 328046 471250 328102
rect 471306 328046 471374 328102
rect 471430 328046 471498 328102
rect 471554 328046 471622 328102
rect 471678 328046 489250 328102
rect 489306 328046 489374 328102
rect 489430 328046 489498 328102
rect 489554 328046 489622 328102
rect 489678 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 64518 327978
rect 64574 327922 64642 327978
rect 64698 327922 95238 327978
rect 95294 327922 95362 327978
rect 95418 327922 125958 327978
rect 126014 327922 126082 327978
rect 126138 327922 156678 327978
rect 156734 327922 156802 327978
rect 156858 327922 187398 327978
rect 187454 327922 187522 327978
rect 187578 327922 218118 327978
rect 218174 327922 218242 327978
rect 218298 327922 248838 327978
rect 248894 327922 248962 327978
rect 249018 327922 279558 327978
rect 279614 327922 279682 327978
rect 279738 327922 310278 327978
rect 310334 327922 310402 327978
rect 310458 327922 340998 327978
rect 341054 327922 341122 327978
rect 341178 327922 363250 327978
rect 363306 327922 363374 327978
rect 363430 327922 363498 327978
rect 363554 327922 363622 327978
rect 363678 327922 371718 327978
rect 371774 327922 371842 327978
rect 371898 327922 381250 327978
rect 381306 327922 381374 327978
rect 381430 327922 381498 327978
rect 381554 327922 381622 327978
rect 381678 327922 399250 327978
rect 399306 327922 399374 327978
rect 399430 327922 399498 327978
rect 399554 327922 399622 327978
rect 399678 327922 402438 327978
rect 402494 327922 402562 327978
rect 402618 327922 433158 327978
rect 433214 327922 433282 327978
rect 433338 327922 435250 327978
rect 435306 327922 435374 327978
rect 435430 327922 435498 327978
rect 435554 327922 435622 327978
rect 435678 327922 453250 327978
rect 453306 327922 453374 327978
rect 453430 327922 453498 327978
rect 453554 327922 453622 327978
rect 453678 327922 471250 327978
rect 471306 327922 471374 327978
rect 471430 327922 471498 327978
rect 471554 327922 471622 327978
rect 471678 327922 489250 327978
rect 489306 327922 489374 327978
rect 489430 327922 489498 327978
rect 489554 327922 489622 327978
rect 489678 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 79878 316350
rect 79934 316294 80002 316350
rect 80058 316294 110598 316350
rect 110654 316294 110722 316350
rect 110778 316294 141318 316350
rect 141374 316294 141442 316350
rect 141498 316294 172038 316350
rect 172094 316294 172162 316350
rect 172218 316294 202758 316350
rect 202814 316294 202882 316350
rect 202938 316294 233478 316350
rect 233534 316294 233602 316350
rect 233658 316294 264198 316350
rect 264254 316294 264322 316350
rect 264378 316294 294918 316350
rect 294974 316294 295042 316350
rect 295098 316294 325638 316350
rect 325694 316294 325762 316350
rect 325818 316294 348970 316350
rect 349026 316294 349094 316350
rect 349150 316294 349218 316350
rect 349274 316294 349342 316350
rect 349398 316294 356358 316350
rect 356414 316294 356482 316350
rect 356538 316294 366970 316350
rect 367026 316294 367094 316350
rect 367150 316294 367218 316350
rect 367274 316294 367342 316350
rect 367398 316294 384970 316350
rect 385026 316294 385094 316350
rect 385150 316294 385218 316350
rect 385274 316294 385342 316350
rect 385398 316294 387078 316350
rect 387134 316294 387202 316350
rect 387258 316294 402970 316350
rect 403026 316294 403094 316350
rect 403150 316294 403218 316350
rect 403274 316294 403342 316350
rect 403398 316294 417798 316350
rect 417854 316294 417922 316350
rect 417978 316294 420970 316350
rect 421026 316294 421094 316350
rect 421150 316294 421218 316350
rect 421274 316294 421342 316350
rect 421398 316294 438970 316350
rect 439026 316294 439094 316350
rect 439150 316294 439218 316350
rect 439274 316294 439342 316350
rect 439398 316294 456970 316350
rect 457026 316294 457094 316350
rect 457150 316294 457218 316350
rect 457274 316294 457342 316350
rect 457398 316294 474970 316350
rect 475026 316294 475094 316350
rect 475150 316294 475218 316350
rect 475274 316294 475342 316350
rect 475398 316294 492970 316350
rect 493026 316294 493094 316350
rect 493150 316294 493218 316350
rect 493274 316294 493342 316350
rect 493398 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 79878 316226
rect 79934 316170 80002 316226
rect 80058 316170 110598 316226
rect 110654 316170 110722 316226
rect 110778 316170 141318 316226
rect 141374 316170 141442 316226
rect 141498 316170 172038 316226
rect 172094 316170 172162 316226
rect 172218 316170 202758 316226
rect 202814 316170 202882 316226
rect 202938 316170 233478 316226
rect 233534 316170 233602 316226
rect 233658 316170 264198 316226
rect 264254 316170 264322 316226
rect 264378 316170 294918 316226
rect 294974 316170 295042 316226
rect 295098 316170 325638 316226
rect 325694 316170 325762 316226
rect 325818 316170 348970 316226
rect 349026 316170 349094 316226
rect 349150 316170 349218 316226
rect 349274 316170 349342 316226
rect 349398 316170 356358 316226
rect 356414 316170 356482 316226
rect 356538 316170 366970 316226
rect 367026 316170 367094 316226
rect 367150 316170 367218 316226
rect 367274 316170 367342 316226
rect 367398 316170 384970 316226
rect 385026 316170 385094 316226
rect 385150 316170 385218 316226
rect 385274 316170 385342 316226
rect 385398 316170 387078 316226
rect 387134 316170 387202 316226
rect 387258 316170 402970 316226
rect 403026 316170 403094 316226
rect 403150 316170 403218 316226
rect 403274 316170 403342 316226
rect 403398 316170 417798 316226
rect 417854 316170 417922 316226
rect 417978 316170 420970 316226
rect 421026 316170 421094 316226
rect 421150 316170 421218 316226
rect 421274 316170 421342 316226
rect 421398 316170 438970 316226
rect 439026 316170 439094 316226
rect 439150 316170 439218 316226
rect 439274 316170 439342 316226
rect 439398 316170 456970 316226
rect 457026 316170 457094 316226
rect 457150 316170 457218 316226
rect 457274 316170 457342 316226
rect 457398 316170 474970 316226
rect 475026 316170 475094 316226
rect 475150 316170 475218 316226
rect 475274 316170 475342 316226
rect 475398 316170 492970 316226
rect 493026 316170 493094 316226
rect 493150 316170 493218 316226
rect 493274 316170 493342 316226
rect 493398 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 79878 316102
rect 79934 316046 80002 316102
rect 80058 316046 110598 316102
rect 110654 316046 110722 316102
rect 110778 316046 141318 316102
rect 141374 316046 141442 316102
rect 141498 316046 172038 316102
rect 172094 316046 172162 316102
rect 172218 316046 202758 316102
rect 202814 316046 202882 316102
rect 202938 316046 233478 316102
rect 233534 316046 233602 316102
rect 233658 316046 264198 316102
rect 264254 316046 264322 316102
rect 264378 316046 294918 316102
rect 294974 316046 295042 316102
rect 295098 316046 325638 316102
rect 325694 316046 325762 316102
rect 325818 316046 348970 316102
rect 349026 316046 349094 316102
rect 349150 316046 349218 316102
rect 349274 316046 349342 316102
rect 349398 316046 356358 316102
rect 356414 316046 356482 316102
rect 356538 316046 366970 316102
rect 367026 316046 367094 316102
rect 367150 316046 367218 316102
rect 367274 316046 367342 316102
rect 367398 316046 384970 316102
rect 385026 316046 385094 316102
rect 385150 316046 385218 316102
rect 385274 316046 385342 316102
rect 385398 316046 387078 316102
rect 387134 316046 387202 316102
rect 387258 316046 402970 316102
rect 403026 316046 403094 316102
rect 403150 316046 403218 316102
rect 403274 316046 403342 316102
rect 403398 316046 417798 316102
rect 417854 316046 417922 316102
rect 417978 316046 420970 316102
rect 421026 316046 421094 316102
rect 421150 316046 421218 316102
rect 421274 316046 421342 316102
rect 421398 316046 438970 316102
rect 439026 316046 439094 316102
rect 439150 316046 439218 316102
rect 439274 316046 439342 316102
rect 439398 316046 456970 316102
rect 457026 316046 457094 316102
rect 457150 316046 457218 316102
rect 457274 316046 457342 316102
rect 457398 316046 474970 316102
rect 475026 316046 475094 316102
rect 475150 316046 475218 316102
rect 475274 316046 475342 316102
rect 475398 316046 492970 316102
rect 493026 316046 493094 316102
rect 493150 316046 493218 316102
rect 493274 316046 493342 316102
rect 493398 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 79878 315978
rect 79934 315922 80002 315978
rect 80058 315922 110598 315978
rect 110654 315922 110722 315978
rect 110778 315922 141318 315978
rect 141374 315922 141442 315978
rect 141498 315922 172038 315978
rect 172094 315922 172162 315978
rect 172218 315922 202758 315978
rect 202814 315922 202882 315978
rect 202938 315922 233478 315978
rect 233534 315922 233602 315978
rect 233658 315922 264198 315978
rect 264254 315922 264322 315978
rect 264378 315922 294918 315978
rect 294974 315922 295042 315978
rect 295098 315922 325638 315978
rect 325694 315922 325762 315978
rect 325818 315922 348970 315978
rect 349026 315922 349094 315978
rect 349150 315922 349218 315978
rect 349274 315922 349342 315978
rect 349398 315922 356358 315978
rect 356414 315922 356482 315978
rect 356538 315922 366970 315978
rect 367026 315922 367094 315978
rect 367150 315922 367218 315978
rect 367274 315922 367342 315978
rect 367398 315922 384970 315978
rect 385026 315922 385094 315978
rect 385150 315922 385218 315978
rect 385274 315922 385342 315978
rect 385398 315922 387078 315978
rect 387134 315922 387202 315978
rect 387258 315922 402970 315978
rect 403026 315922 403094 315978
rect 403150 315922 403218 315978
rect 403274 315922 403342 315978
rect 403398 315922 417798 315978
rect 417854 315922 417922 315978
rect 417978 315922 420970 315978
rect 421026 315922 421094 315978
rect 421150 315922 421218 315978
rect 421274 315922 421342 315978
rect 421398 315922 438970 315978
rect 439026 315922 439094 315978
rect 439150 315922 439218 315978
rect 439274 315922 439342 315978
rect 439398 315922 456970 315978
rect 457026 315922 457094 315978
rect 457150 315922 457218 315978
rect 457274 315922 457342 315978
rect 457398 315922 474970 315978
rect 475026 315922 475094 315978
rect 475150 315922 475218 315978
rect 475274 315922 475342 315978
rect 475398 315922 492970 315978
rect 493026 315922 493094 315978
rect 493150 315922 493218 315978
rect 493274 315922 493342 315978
rect 493398 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 64518 310350
rect 64574 310294 64642 310350
rect 64698 310294 95238 310350
rect 95294 310294 95362 310350
rect 95418 310294 125958 310350
rect 126014 310294 126082 310350
rect 126138 310294 156678 310350
rect 156734 310294 156802 310350
rect 156858 310294 187398 310350
rect 187454 310294 187522 310350
rect 187578 310294 218118 310350
rect 218174 310294 218242 310350
rect 218298 310294 248838 310350
rect 248894 310294 248962 310350
rect 249018 310294 279558 310350
rect 279614 310294 279682 310350
rect 279738 310294 310278 310350
rect 310334 310294 310402 310350
rect 310458 310294 340998 310350
rect 341054 310294 341122 310350
rect 341178 310294 363250 310350
rect 363306 310294 363374 310350
rect 363430 310294 363498 310350
rect 363554 310294 363622 310350
rect 363678 310294 371718 310350
rect 371774 310294 371842 310350
rect 371898 310294 381250 310350
rect 381306 310294 381374 310350
rect 381430 310294 381498 310350
rect 381554 310294 381622 310350
rect 381678 310294 399250 310350
rect 399306 310294 399374 310350
rect 399430 310294 399498 310350
rect 399554 310294 399622 310350
rect 399678 310294 402438 310350
rect 402494 310294 402562 310350
rect 402618 310294 433158 310350
rect 433214 310294 433282 310350
rect 433338 310294 435250 310350
rect 435306 310294 435374 310350
rect 435430 310294 435498 310350
rect 435554 310294 435622 310350
rect 435678 310294 453250 310350
rect 453306 310294 453374 310350
rect 453430 310294 453498 310350
rect 453554 310294 453622 310350
rect 453678 310294 471250 310350
rect 471306 310294 471374 310350
rect 471430 310294 471498 310350
rect 471554 310294 471622 310350
rect 471678 310294 489250 310350
rect 489306 310294 489374 310350
rect 489430 310294 489498 310350
rect 489554 310294 489622 310350
rect 489678 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 64518 310226
rect 64574 310170 64642 310226
rect 64698 310170 95238 310226
rect 95294 310170 95362 310226
rect 95418 310170 125958 310226
rect 126014 310170 126082 310226
rect 126138 310170 156678 310226
rect 156734 310170 156802 310226
rect 156858 310170 187398 310226
rect 187454 310170 187522 310226
rect 187578 310170 218118 310226
rect 218174 310170 218242 310226
rect 218298 310170 248838 310226
rect 248894 310170 248962 310226
rect 249018 310170 279558 310226
rect 279614 310170 279682 310226
rect 279738 310170 310278 310226
rect 310334 310170 310402 310226
rect 310458 310170 340998 310226
rect 341054 310170 341122 310226
rect 341178 310170 363250 310226
rect 363306 310170 363374 310226
rect 363430 310170 363498 310226
rect 363554 310170 363622 310226
rect 363678 310170 371718 310226
rect 371774 310170 371842 310226
rect 371898 310170 381250 310226
rect 381306 310170 381374 310226
rect 381430 310170 381498 310226
rect 381554 310170 381622 310226
rect 381678 310170 399250 310226
rect 399306 310170 399374 310226
rect 399430 310170 399498 310226
rect 399554 310170 399622 310226
rect 399678 310170 402438 310226
rect 402494 310170 402562 310226
rect 402618 310170 433158 310226
rect 433214 310170 433282 310226
rect 433338 310170 435250 310226
rect 435306 310170 435374 310226
rect 435430 310170 435498 310226
rect 435554 310170 435622 310226
rect 435678 310170 453250 310226
rect 453306 310170 453374 310226
rect 453430 310170 453498 310226
rect 453554 310170 453622 310226
rect 453678 310170 471250 310226
rect 471306 310170 471374 310226
rect 471430 310170 471498 310226
rect 471554 310170 471622 310226
rect 471678 310170 489250 310226
rect 489306 310170 489374 310226
rect 489430 310170 489498 310226
rect 489554 310170 489622 310226
rect 489678 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 64518 310102
rect 64574 310046 64642 310102
rect 64698 310046 95238 310102
rect 95294 310046 95362 310102
rect 95418 310046 125958 310102
rect 126014 310046 126082 310102
rect 126138 310046 156678 310102
rect 156734 310046 156802 310102
rect 156858 310046 187398 310102
rect 187454 310046 187522 310102
rect 187578 310046 218118 310102
rect 218174 310046 218242 310102
rect 218298 310046 248838 310102
rect 248894 310046 248962 310102
rect 249018 310046 279558 310102
rect 279614 310046 279682 310102
rect 279738 310046 310278 310102
rect 310334 310046 310402 310102
rect 310458 310046 340998 310102
rect 341054 310046 341122 310102
rect 341178 310046 363250 310102
rect 363306 310046 363374 310102
rect 363430 310046 363498 310102
rect 363554 310046 363622 310102
rect 363678 310046 371718 310102
rect 371774 310046 371842 310102
rect 371898 310046 381250 310102
rect 381306 310046 381374 310102
rect 381430 310046 381498 310102
rect 381554 310046 381622 310102
rect 381678 310046 399250 310102
rect 399306 310046 399374 310102
rect 399430 310046 399498 310102
rect 399554 310046 399622 310102
rect 399678 310046 402438 310102
rect 402494 310046 402562 310102
rect 402618 310046 433158 310102
rect 433214 310046 433282 310102
rect 433338 310046 435250 310102
rect 435306 310046 435374 310102
rect 435430 310046 435498 310102
rect 435554 310046 435622 310102
rect 435678 310046 453250 310102
rect 453306 310046 453374 310102
rect 453430 310046 453498 310102
rect 453554 310046 453622 310102
rect 453678 310046 471250 310102
rect 471306 310046 471374 310102
rect 471430 310046 471498 310102
rect 471554 310046 471622 310102
rect 471678 310046 489250 310102
rect 489306 310046 489374 310102
rect 489430 310046 489498 310102
rect 489554 310046 489622 310102
rect 489678 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 64518 309978
rect 64574 309922 64642 309978
rect 64698 309922 95238 309978
rect 95294 309922 95362 309978
rect 95418 309922 125958 309978
rect 126014 309922 126082 309978
rect 126138 309922 156678 309978
rect 156734 309922 156802 309978
rect 156858 309922 187398 309978
rect 187454 309922 187522 309978
rect 187578 309922 218118 309978
rect 218174 309922 218242 309978
rect 218298 309922 248838 309978
rect 248894 309922 248962 309978
rect 249018 309922 279558 309978
rect 279614 309922 279682 309978
rect 279738 309922 310278 309978
rect 310334 309922 310402 309978
rect 310458 309922 340998 309978
rect 341054 309922 341122 309978
rect 341178 309922 363250 309978
rect 363306 309922 363374 309978
rect 363430 309922 363498 309978
rect 363554 309922 363622 309978
rect 363678 309922 371718 309978
rect 371774 309922 371842 309978
rect 371898 309922 381250 309978
rect 381306 309922 381374 309978
rect 381430 309922 381498 309978
rect 381554 309922 381622 309978
rect 381678 309922 399250 309978
rect 399306 309922 399374 309978
rect 399430 309922 399498 309978
rect 399554 309922 399622 309978
rect 399678 309922 402438 309978
rect 402494 309922 402562 309978
rect 402618 309922 433158 309978
rect 433214 309922 433282 309978
rect 433338 309922 435250 309978
rect 435306 309922 435374 309978
rect 435430 309922 435498 309978
rect 435554 309922 435622 309978
rect 435678 309922 453250 309978
rect 453306 309922 453374 309978
rect 453430 309922 453498 309978
rect 453554 309922 453622 309978
rect 453678 309922 471250 309978
rect 471306 309922 471374 309978
rect 471430 309922 471498 309978
rect 471554 309922 471622 309978
rect 471678 309922 489250 309978
rect 489306 309922 489374 309978
rect 489430 309922 489498 309978
rect 489554 309922 489622 309978
rect 489678 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 79878 298350
rect 79934 298294 80002 298350
rect 80058 298294 110598 298350
rect 110654 298294 110722 298350
rect 110778 298294 141318 298350
rect 141374 298294 141442 298350
rect 141498 298294 172038 298350
rect 172094 298294 172162 298350
rect 172218 298294 202758 298350
rect 202814 298294 202882 298350
rect 202938 298294 233478 298350
rect 233534 298294 233602 298350
rect 233658 298294 264198 298350
rect 264254 298294 264322 298350
rect 264378 298294 294918 298350
rect 294974 298294 295042 298350
rect 295098 298294 325638 298350
rect 325694 298294 325762 298350
rect 325818 298294 348970 298350
rect 349026 298294 349094 298350
rect 349150 298294 349218 298350
rect 349274 298294 349342 298350
rect 349398 298294 356358 298350
rect 356414 298294 356482 298350
rect 356538 298294 366970 298350
rect 367026 298294 367094 298350
rect 367150 298294 367218 298350
rect 367274 298294 367342 298350
rect 367398 298294 384970 298350
rect 385026 298294 385094 298350
rect 385150 298294 385218 298350
rect 385274 298294 385342 298350
rect 385398 298294 387078 298350
rect 387134 298294 387202 298350
rect 387258 298294 402970 298350
rect 403026 298294 403094 298350
rect 403150 298294 403218 298350
rect 403274 298294 403342 298350
rect 403398 298294 417798 298350
rect 417854 298294 417922 298350
rect 417978 298294 420970 298350
rect 421026 298294 421094 298350
rect 421150 298294 421218 298350
rect 421274 298294 421342 298350
rect 421398 298294 438970 298350
rect 439026 298294 439094 298350
rect 439150 298294 439218 298350
rect 439274 298294 439342 298350
rect 439398 298294 456970 298350
rect 457026 298294 457094 298350
rect 457150 298294 457218 298350
rect 457274 298294 457342 298350
rect 457398 298294 474970 298350
rect 475026 298294 475094 298350
rect 475150 298294 475218 298350
rect 475274 298294 475342 298350
rect 475398 298294 492970 298350
rect 493026 298294 493094 298350
rect 493150 298294 493218 298350
rect 493274 298294 493342 298350
rect 493398 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 79878 298226
rect 79934 298170 80002 298226
rect 80058 298170 110598 298226
rect 110654 298170 110722 298226
rect 110778 298170 141318 298226
rect 141374 298170 141442 298226
rect 141498 298170 172038 298226
rect 172094 298170 172162 298226
rect 172218 298170 202758 298226
rect 202814 298170 202882 298226
rect 202938 298170 233478 298226
rect 233534 298170 233602 298226
rect 233658 298170 264198 298226
rect 264254 298170 264322 298226
rect 264378 298170 294918 298226
rect 294974 298170 295042 298226
rect 295098 298170 325638 298226
rect 325694 298170 325762 298226
rect 325818 298170 348970 298226
rect 349026 298170 349094 298226
rect 349150 298170 349218 298226
rect 349274 298170 349342 298226
rect 349398 298170 356358 298226
rect 356414 298170 356482 298226
rect 356538 298170 366970 298226
rect 367026 298170 367094 298226
rect 367150 298170 367218 298226
rect 367274 298170 367342 298226
rect 367398 298170 384970 298226
rect 385026 298170 385094 298226
rect 385150 298170 385218 298226
rect 385274 298170 385342 298226
rect 385398 298170 387078 298226
rect 387134 298170 387202 298226
rect 387258 298170 402970 298226
rect 403026 298170 403094 298226
rect 403150 298170 403218 298226
rect 403274 298170 403342 298226
rect 403398 298170 417798 298226
rect 417854 298170 417922 298226
rect 417978 298170 420970 298226
rect 421026 298170 421094 298226
rect 421150 298170 421218 298226
rect 421274 298170 421342 298226
rect 421398 298170 438970 298226
rect 439026 298170 439094 298226
rect 439150 298170 439218 298226
rect 439274 298170 439342 298226
rect 439398 298170 456970 298226
rect 457026 298170 457094 298226
rect 457150 298170 457218 298226
rect 457274 298170 457342 298226
rect 457398 298170 474970 298226
rect 475026 298170 475094 298226
rect 475150 298170 475218 298226
rect 475274 298170 475342 298226
rect 475398 298170 492970 298226
rect 493026 298170 493094 298226
rect 493150 298170 493218 298226
rect 493274 298170 493342 298226
rect 493398 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 79878 298102
rect 79934 298046 80002 298102
rect 80058 298046 110598 298102
rect 110654 298046 110722 298102
rect 110778 298046 141318 298102
rect 141374 298046 141442 298102
rect 141498 298046 172038 298102
rect 172094 298046 172162 298102
rect 172218 298046 202758 298102
rect 202814 298046 202882 298102
rect 202938 298046 233478 298102
rect 233534 298046 233602 298102
rect 233658 298046 264198 298102
rect 264254 298046 264322 298102
rect 264378 298046 294918 298102
rect 294974 298046 295042 298102
rect 295098 298046 325638 298102
rect 325694 298046 325762 298102
rect 325818 298046 348970 298102
rect 349026 298046 349094 298102
rect 349150 298046 349218 298102
rect 349274 298046 349342 298102
rect 349398 298046 356358 298102
rect 356414 298046 356482 298102
rect 356538 298046 366970 298102
rect 367026 298046 367094 298102
rect 367150 298046 367218 298102
rect 367274 298046 367342 298102
rect 367398 298046 384970 298102
rect 385026 298046 385094 298102
rect 385150 298046 385218 298102
rect 385274 298046 385342 298102
rect 385398 298046 387078 298102
rect 387134 298046 387202 298102
rect 387258 298046 402970 298102
rect 403026 298046 403094 298102
rect 403150 298046 403218 298102
rect 403274 298046 403342 298102
rect 403398 298046 417798 298102
rect 417854 298046 417922 298102
rect 417978 298046 420970 298102
rect 421026 298046 421094 298102
rect 421150 298046 421218 298102
rect 421274 298046 421342 298102
rect 421398 298046 438970 298102
rect 439026 298046 439094 298102
rect 439150 298046 439218 298102
rect 439274 298046 439342 298102
rect 439398 298046 456970 298102
rect 457026 298046 457094 298102
rect 457150 298046 457218 298102
rect 457274 298046 457342 298102
rect 457398 298046 474970 298102
rect 475026 298046 475094 298102
rect 475150 298046 475218 298102
rect 475274 298046 475342 298102
rect 475398 298046 492970 298102
rect 493026 298046 493094 298102
rect 493150 298046 493218 298102
rect 493274 298046 493342 298102
rect 493398 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 79878 297978
rect 79934 297922 80002 297978
rect 80058 297922 110598 297978
rect 110654 297922 110722 297978
rect 110778 297922 141318 297978
rect 141374 297922 141442 297978
rect 141498 297922 172038 297978
rect 172094 297922 172162 297978
rect 172218 297922 202758 297978
rect 202814 297922 202882 297978
rect 202938 297922 233478 297978
rect 233534 297922 233602 297978
rect 233658 297922 264198 297978
rect 264254 297922 264322 297978
rect 264378 297922 294918 297978
rect 294974 297922 295042 297978
rect 295098 297922 325638 297978
rect 325694 297922 325762 297978
rect 325818 297922 348970 297978
rect 349026 297922 349094 297978
rect 349150 297922 349218 297978
rect 349274 297922 349342 297978
rect 349398 297922 356358 297978
rect 356414 297922 356482 297978
rect 356538 297922 366970 297978
rect 367026 297922 367094 297978
rect 367150 297922 367218 297978
rect 367274 297922 367342 297978
rect 367398 297922 384970 297978
rect 385026 297922 385094 297978
rect 385150 297922 385218 297978
rect 385274 297922 385342 297978
rect 385398 297922 387078 297978
rect 387134 297922 387202 297978
rect 387258 297922 402970 297978
rect 403026 297922 403094 297978
rect 403150 297922 403218 297978
rect 403274 297922 403342 297978
rect 403398 297922 417798 297978
rect 417854 297922 417922 297978
rect 417978 297922 420970 297978
rect 421026 297922 421094 297978
rect 421150 297922 421218 297978
rect 421274 297922 421342 297978
rect 421398 297922 438970 297978
rect 439026 297922 439094 297978
rect 439150 297922 439218 297978
rect 439274 297922 439342 297978
rect 439398 297922 456970 297978
rect 457026 297922 457094 297978
rect 457150 297922 457218 297978
rect 457274 297922 457342 297978
rect 457398 297922 474970 297978
rect 475026 297922 475094 297978
rect 475150 297922 475218 297978
rect 475274 297922 475342 297978
rect 475398 297922 492970 297978
rect 493026 297922 493094 297978
rect 493150 297922 493218 297978
rect 493274 297922 493342 297978
rect 493398 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 64518 292350
rect 64574 292294 64642 292350
rect 64698 292294 95238 292350
rect 95294 292294 95362 292350
rect 95418 292294 125958 292350
rect 126014 292294 126082 292350
rect 126138 292294 156678 292350
rect 156734 292294 156802 292350
rect 156858 292294 187398 292350
rect 187454 292294 187522 292350
rect 187578 292294 218118 292350
rect 218174 292294 218242 292350
rect 218298 292294 248838 292350
rect 248894 292294 248962 292350
rect 249018 292294 279558 292350
rect 279614 292294 279682 292350
rect 279738 292294 310278 292350
rect 310334 292294 310402 292350
rect 310458 292294 340998 292350
rect 341054 292294 341122 292350
rect 341178 292294 363250 292350
rect 363306 292294 363374 292350
rect 363430 292294 363498 292350
rect 363554 292294 363622 292350
rect 363678 292294 371718 292350
rect 371774 292294 371842 292350
rect 371898 292294 381250 292350
rect 381306 292294 381374 292350
rect 381430 292294 381498 292350
rect 381554 292294 381622 292350
rect 381678 292294 399250 292350
rect 399306 292294 399374 292350
rect 399430 292294 399498 292350
rect 399554 292294 399622 292350
rect 399678 292294 402438 292350
rect 402494 292294 402562 292350
rect 402618 292294 433158 292350
rect 433214 292294 433282 292350
rect 433338 292294 435250 292350
rect 435306 292294 435374 292350
rect 435430 292294 435498 292350
rect 435554 292294 435622 292350
rect 435678 292294 453250 292350
rect 453306 292294 453374 292350
rect 453430 292294 453498 292350
rect 453554 292294 453622 292350
rect 453678 292294 471250 292350
rect 471306 292294 471374 292350
rect 471430 292294 471498 292350
rect 471554 292294 471622 292350
rect 471678 292294 489250 292350
rect 489306 292294 489374 292350
rect 489430 292294 489498 292350
rect 489554 292294 489622 292350
rect 489678 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 64518 292226
rect 64574 292170 64642 292226
rect 64698 292170 95238 292226
rect 95294 292170 95362 292226
rect 95418 292170 125958 292226
rect 126014 292170 126082 292226
rect 126138 292170 156678 292226
rect 156734 292170 156802 292226
rect 156858 292170 187398 292226
rect 187454 292170 187522 292226
rect 187578 292170 218118 292226
rect 218174 292170 218242 292226
rect 218298 292170 248838 292226
rect 248894 292170 248962 292226
rect 249018 292170 279558 292226
rect 279614 292170 279682 292226
rect 279738 292170 310278 292226
rect 310334 292170 310402 292226
rect 310458 292170 340998 292226
rect 341054 292170 341122 292226
rect 341178 292170 363250 292226
rect 363306 292170 363374 292226
rect 363430 292170 363498 292226
rect 363554 292170 363622 292226
rect 363678 292170 371718 292226
rect 371774 292170 371842 292226
rect 371898 292170 381250 292226
rect 381306 292170 381374 292226
rect 381430 292170 381498 292226
rect 381554 292170 381622 292226
rect 381678 292170 399250 292226
rect 399306 292170 399374 292226
rect 399430 292170 399498 292226
rect 399554 292170 399622 292226
rect 399678 292170 402438 292226
rect 402494 292170 402562 292226
rect 402618 292170 433158 292226
rect 433214 292170 433282 292226
rect 433338 292170 435250 292226
rect 435306 292170 435374 292226
rect 435430 292170 435498 292226
rect 435554 292170 435622 292226
rect 435678 292170 453250 292226
rect 453306 292170 453374 292226
rect 453430 292170 453498 292226
rect 453554 292170 453622 292226
rect 453678 292170 471250 292226
rect 471306 292170 471374 292226
rect 471430 292170 471498 292226
rect 471554 292170 471622 292226
rect 471678 292170 489250 292226
rect 489306 292170 489374 292226
rect 489430 292170 489498 292226
rect 489554 292170 489622 292226
rect 489678 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 64518 292102
rect 64574 292046 64642 292102
rect 64698 292046 95238 292102
rect 95294 292046 95362 292102
rect 95418 292046 125958 292102
rect 126014 292046 126082 292102
rect 126138 292046 156678 292102
rect 156734 292046 156802 292102
rect 156858 292046 187398 292102
rect 187454 292046 187522 292102
rect 187578 292046 218118 292102
rect 218174 292046 218242 292102
rect 218298 292046 248838 292102
rect 248894 292046 248962 292102
rect 249018 292046 279558 292102
rect 279614 292046 279682 292102
rect 279738 292046 310278 292102
rect 310334 292046 310402 292102
rect 310458 292046 340998 292102
rect 341054 292046 341122 292102
rect 341178 292046 363250 292102
rect 363306 292046 363374 292102
rect 363430 292046 363498 292102
rect 363554 292046 363622 292102
rect 363678 292046 371718 292102
rect 371774 292046 371842 292102
rect 371898 292046 381250 292102
rect 381306 292046 381374 292102
rect 381430 292046 381498 292102
rect 381554 292046 381622 292102
rect 381678 292046 399250 292102
rect 399306 292046 399374 292102
rect 399430 292046 399498 292102
rect 399554 292046 399622 292102
rect 399678 292046 402438 292102
rect 402494 292046 402562 292102
rect 402618 292046 433158 292102
rect 433214 292046 433282 292102
rect 433338 292046 435250 292102
rect 435306 292046 435374 292102
rect 435430 292046 435498 292102
rect 435554 292046 435622 292102
rect 435678 292046 453250 292102
rect 453306 292046 453374 292102
rect 453430 292046 453498 292102
rect 453554 292046 453622 292102
rect 453678 292046 471250 292102
rect 471306 292046 471374 292102
rect 471430 292046 471498 292102
rect 471554 292046 471622 292102
rect 471678 292046 489250 292102
rect 489306 292046 489374 292102
rect 489430 292046 489498 292102
rect 489554 292046 489622 292102
rect 489678 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 64518 291978
rect 64574 291922 64642 291978
rect 64698 291922 95238 291978
rect 95294 291922 95362 291978
rect 95418 291922 125958 291978
rect 126014 291922 126082 291978
rect 126138 291922 156678 291978
rect 156734 291922 156802 291978
rect 156858 291922 187398 291978
rect 187454 291922 187522 291978
rect 187578 291922 218118 291978
rect 218174 291922 218242 291978
rect 218298 291922 248838 291978
rect 248894 291922 248962 291978
rect 249018 291922 279558 291978
rect 279614 291922 279682 291978
rect 279738 291922 310278 291978
rect 310334 291922 310402 291978
rect 310458 291922 340998 291978
rect 341054 291922 341122 291978
rect 341178 291922 363250 291978
rect 363306 291922 363374 291978
rect 363430 291922 363498 291978
rect 363554 291922 363622 291978
rect 363678 291922 371718 291978
rect 371774 291922 371842 291978
rect 371898 291922 381250 291978
rect 381306 291922 381374 291978
rect 381430 291922 381498 291978
rect 381554 291922 381622 291978
rect 381678 291922 399250 291978
rect 399306 291922 399374 291978
rect 399430 291922 399498 291978
rect 399554 291922 399622 291978
rect 399678 291922 402438 291978
rect 402494 291922 402562 291978
rect 402618 291922 433158 291978
rect 433214 291922 433282 291978
rect 433338 291922 435250 291978
rect 435306 291922 435374 291978
rect 435430 291922 435498 291978
rect 435554 291922 435622 291978
rect 435678 291922 453250 291978
rect 453306 291922 453374 291978
rect 453430 291922 453498 291978
rect 453554 291922 453622 291978
rect 453678 291922 471250 291978
rect 471306 291922 471374 291978
rect 471430 291922 471498 291978
rect 471554 291922 471622 291978
rect 471678 291922 489250 291978
rect 489306 291922 489374 291978
rect 489430 291922 489498 291978
rect 489554 291922 489622 291978
rect 489678 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 79878 280350
rect 79934 280294 80002 280350
rect 80058 280294 110598 280350
rect 110654 280294 110722 280350
rect 110778 280294 141318 280350
rect 141374 280294 141442 280350
rect 141498 280294 172038 280350
rect 172094 280294 172162 280350
rect 172218 280294 202758 280350
rect 202814 280294 202882 280350
rect 202938 280294 233478 280350
rect 233534 280294 233602 280350
rect 233658 280294 264198 280350
rect 264254 280294 264322 280350
rect 264378 280294 294918 280350
rect 294974 280294 295042 280350
rect 295098 280294 325638 280350
rect 325694 280294 325762 280350
rect 325818 280294 348970 280350
rect 349026 280294 349094 280350
rect 349150 280294 349218 280350
rect 349274 280294 349342 280350
rect 349398 280294 356358 280350
rect 356414 280294 356482 280350
rect 356538 280294 366970 280350
rect 367026 280294 367094 280350
rect 367150 280294 367218 280350
rect 367274 280294 367342 280350
rect 367398 280294 384970 280350
rect 385026 280294 385094 280350
rect 385150 280294 385218 280350
rect 385274 280294 385342 280350
rect 385398 280294 387078 280350
rect 387134 280294 387202 280350
rect 387258 280294 402970 280350
rect 403026 280294 403094 280350
rect 403150 280294 403218 280350
rect 403274 280294 403342 280350
rect 403398 280294 417798 280350
rect 417854 280294 417922 280350
rect 417978 280294 420970 280350
rect 421026 280294 421094 280350
rect 421150 280294 421218 280350
rect 421274 280294 421342 280350
rect 421398 280294 438970 280350
rect 439026 280294 439094 280350
rect 439150 280294 439218 280350
rect 439274 280294 439342 280350
rect 439398 280294 456970 280350
rect 457026 280294 457094 280350
rect 457150 280294 457218 280350
rect 457274 280294 457342 280350
rect 457398 280294 474970 280350
rect 475026 280294 475094 280350
rect 475150 280294 475218 280350
rect 475274 280294 475342 280350
rect 475398 280294 492970 280350
rect 493026 280294 493094 280350
rect 493150 280294 493218 280350
rect 493274 280294 493342 280350
rect 493398 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 79878 280226
rect 79934 280170 80002 280226
rect 80058 280170 110598 280226
rect 110654 280170 110722 280226
rect 110778 280170 141318 280226
rect 141374 280170 141442 280226
rect 141498 280170 172038 280226
rect 172094 280170 172162 280226
rect 172218 280170 202758 280226
rect 202814 280170 202882 280226
rect 202938 280170 233478 280226
rect 233534 280170 233602 280226
rect 233658 280170 264198 280226
rect 264254 280170 264322 280226
rect 264378 280170 294918 280226
rect 294974 280170 295042 280226
rect 295098 280170 325638 280226
rect 325694 280170 325762 280226
rect 325818 280170 348970 280226
rect 349026 280170 349094 280226
rect 349150 280170 349218 280226
rect 349274 280170 349342 280226
rect 349398 280170 356358 280226
rect 356414 280170 356482 280226
rect 356538 280170 366970 280226
rect 367026 280170 367094 280226
rect 367150 280170 367218 280226
rect 367274 280170 367342 280226
rect 367398 280170 384970 280226
rect 385026 280170 385094 280226
rect 385150 280170 385218 280226
rect 385274 280170 385342 280226
rect 385398 280170 387078 280226
rect 387134 280170 387202 280226
rect 387258 280170 402970 280226
rect 403026 280170 403094 280226
rect 403150 280170 403218 280226
rect 403274 280170 403342 280226
rect 403398 280170 417798 280226
rect 417854 280170 417922 280226
rect 417978 280170 420970 280226
rect 421026 280170 421094 280226
rect 421150 280170 421218 280226
rect 421274 280170 421342 280226
rect 421398 280170 438970 280226
rect 439026 280170 439094 280226
rect 439150 280170 439218 280226
rect 439274 280170 439342 280226
rect 439398 280170 456970 280226
rect 457026 280170 457094 280226
rect 457150 280170 457218 280226
rect 457274 280170 457342 280226
rect 457398 280170 474970 280226
rect 475026 280170 475094 280226
rect 475150 280170 475218 280226
rect 475274 280170 475342 280226
rect 475398 280170 492970 280226
rect 493026 280170 493094 280226
rect 493150 280170 493218 280226
rect 493274 280170 493342 280226
rect 493398 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 79878 280102
rect 79934 280046 80002 280102
rect 80058 280046 110598 280102
rect 110654 280046 110722 280102
rect 110778 280046 141318 280102
rect 141374 280046 141442 280102
rect 141498 280046 172038 280102
rect 172094 280046 172162 280102
rect 172218 280046 202758 280102
rect 202814 280046 202882 280102
rect 202938 280046 233478 280102
rect 233534 280046 233602 280102
rect 233658 280046 264198 280102
rect 264254 280046 264322 280102
rect 264378 280046 294918 280102
rect 294974 280046 295042 280102
rect 295098 280046 325638 280102
rect 325694 280046 325762 280102
rect 325818 280046 348970 280102
rect 349026 280046 349094 280102
rect 349150 280046 349218 280102
rect 349274 280046 349342 280102
rect 349398 280046 356358 280102
rect 356414 280046 356482 280102
rect 356538 280046 366970 280102
rect 367026 280046 367094 280102
rect 367150 280046 367218 280102
rect 367274 280046 367342 280102
rect 367398 280046 384970 280102
rect 385026 280046 385094 280102
rect 385150 280046 385218 280102
rect 385274 280046 385342 280102
rect 385398 280046 387078 280102
rect 387134 280046 387202 280102
rect 387258 280046 402970 280102
rect 403026 280046 403094 280102
rect 403150 280046 403218 280102
rect 403274 280046 403342 280102
rect 403398 280046 417798 280102
rect 417854 280046 417922 280102
rect 417978 280046 420970 280102
rect 421026 280046 421094 280102
rect 421150 280046 421218 280102
rect 421274 280046 421342 280102
rect 421398 280046 438970 280102
rect 439026 280046 439094 280102
rect 439150 280046 439218 280102
rect 439274 280046 439342 280102
rect 439398 280046 456970 280102
rect 457026 280046 457094 280102
rect 457150 280046 457218 280102
rect 457274 280046 457342 280102
rect 457398 280046 474970 280102
rect 475026 280046 475094 280102
rect 475150 280046 475218 280102
rect 475274 280046 475342 280102
rect 475398 280046 492970 280102
rect 493026 280046 493094 280102
rect 493150 280046 493218 280102
rect 493274 280046 493342 280102
rect 493398 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 79878 279978
rect 79934 279922 80002 279978
rect 80058 279922 110598 279978
rect 110654 279922 110722 279978
rect 110778 279922 141318 279978
rect 141374 279922 141442 279978
rect 141498 279922 172038 279978
rect 172094 279922 172162 279978
rect 172218 279922 202758 279978
rect 202814 279922 202882 279978
rect 202938 279922 233478 279978
rect 233534 279922 233602 279978
rect 233658 279922 264198 279978
rect 264254 279922 264322 279978
rect 264378 279922 294918 279978
rect 294974 279922 295042 279978
rect 295098 279922 325638 279978
rect 325694 279922 325762 279978
rect 325818 279922 348970 279978
rect 349026 279922 349094 279978
rect 349150 279922 349218 279978
rect 349274 279922 349342 279978
rect 349398 279922 356358 279978
rect 356414 279922 356482 279978
rect 356538 279922 366970 279978
rect 367026 279922 367094 279978
rect 367150 279922 367218 279978
rect 367274 279922 367342 279978
rect 367398 279922 384970 279978
rect 385026 279922 385094 279978
rect 385150 279922 385218 279978
rect 385274 279922 385342 279978
rect 385398 279922 387078 279978
rect 387134 279922 387202 279978
rect 387258 279922 402970 279978
rect 403026 279922 403094 279978
rect 403150 279922 403218 279978
rect 403274 279922 403342 279978
rect 403398 279922 417798 279978
rect 417854 279922 417922 279978
rect 417978 279922 420970 279978
rect 421026 279922 421094 279978
rect 421150 279922 421218 279978
rect 421274 279922 421342 279978
rect 421398 279922 438970 279978
rect 439026 279922 439094 279978
rect 439150 279922 439218 279978
rect 439274 279922 439342 279978
rect 439398 279922 456970 279978
rect 457026 279922 457094 279978
rect 457150 279922 457218 279978
rect 457274 279922 457342 279978
rect 457398 279922 474970 279978
rect 475026 279922 475094 279978
rect 475150 279922 475218 279978
rect 475274 279922 475342 279978
rect 475398 279922 492970 279978
rect 493026 279922 493094 279978
rect 493150 279922 493218 279978
rect 493274 279922 493342 279978
rect 493398 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 64518 274350
rect 64574 274294 64642 274350
rect 64698 274294 95238 274350
rect 95294 274294 95362 274350
rect 95418 274294 125958 274350
rect 126014 274294 126082 274350
rect 126138 274294 156678 274350
rect 156734 274294 156802 274350
rect 156858 274294 187398 274350
rect 187454 274294 187522 274350
rect 187578 274294 218118 274350
rect 218174 274294 218242 274350
rect 218298 274294 248838 274350
rect 248894 274294 248962 274350
rect 249018 274294 279558 274350
rect 279614 274294 279682 274350
rect 279738 274294 310278 274350
rect 310334 274294 310402 274350
rect 310458 274294 340998 274350
rect 341054 274294 341122 274350
rect 341178 274294 363250 274350
rect 363306 274294 363374 274350
rect 363430 274294 363498 274350
rect 363554 274294 363622 274350
rect 363678 274294 371718 274350
rect 371774 274294 371842 274350
rect 371898 274294 381250 274350
rect 381306 274294 381374 274350
rect 381430 274294 381498 274350
rect 381554 274294 381622 274350
rect 381678 274294 399250 274350
rect 399306 274294 399374 274350
rect 399430 274294 399498 274350
rect 399554 274294 399622 274350
rect 399678 274294 402438 274350
rect 402494 274294 402562 274350
rect 402618 274294 433158 274350
rect 433214 274294 433282 274350
rect 433338 274294 435250 274350
rect 435306 274294 435374 274350
rect 435430 274294 435498 274350
rect 435554 274294 435622 274350
rect 435678 274294 453250 274350
rect 453306 274294 453374 274350
rect 453430 274294 453498 274350
rect 453554 274294 453622 274350
rect 453678 274294 471250 274350
rect 471306 274294 471374 274350
rect 471430 274294 471498 274350
rect 471554 274294 471622 274350
rect 471678 274294 489250 274350
rect 489306 274294 489374 274350
rect 489430 274294 489498 274350
rect 489554 274294 489622 274350
rect 489678 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 64518 274226
rect 64574 274170 64642 274226
rect 64698 274170 95238 274226
rect 95294 274170 95362 274226
rect 95418 274170 125958 274226
rect 126014 274170 126082 274226
rect 126138 274170 156678 274226
rect 156734 274170 156802 274226
rect 156858 274170 187398 274226
rect 187454 274170 187522 274226
rect 187578 274170 218118 274226
rect 218174 274170 218242 274226
rect 218298 274170 248838 274226
rect 248894 274170 248962 274226
rect 249018 274170 279558 274226
rect 279614 274170 279682 274226
rect 279738 274170 310278 274226
rect 310334 274170 310402 274226
rect 310458 274170 340998 274226
rect 341054 274170 341122 274226
rect 341178 274170 363250 274226
rect 363306 274170 363374 274226
rect 363430 274170 363498 274226
rect 363554 274170 363622 274226
rect 363678 274170 371718 274226
rect 371774 274170 371842 274226
rect 371898 274170 381250 274226
rect 381306 274170 381374 274226
rect 381430 274170 381498 274226
rect 381554 274170 381622 274226
rect 381678 274170 399250 274226
rect 399306 274170 399374 274226
rect 399430 274170 399498 274226
rect 399554 274170 399622 274226
rect 399678 274170 402438 274226
rect 402494 274170 402562 274226
rect 402618 274170 433158 274226
rect 433214 274170 433282 274226
rect 433338 274170 435250 274226
rect 435306 274170 435374 274226
rect 435430 274170 435498 274226
rect 435554 274170 435622 274226
rect 435678 274170 453250 274226
rect 453306 274170 453374 274226
rect 453430 274170 453498 274226
rect 453554 274170 453622 274226
rect 453678 274170 471250 274226
rect 471306 274170 471374 274226
rect 471430 274170 471498 274226
rect 471554 274170 471622 274226
rect 471678 274170 489250 274226
rect 489306 274170 489374 274226
rect 489430 274170 489498 274226
rect 489554 274170 489622 274226
rect 489678 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 64518 274102
rect 64574 274046 64642 274102
rect 64698 274046 95238 274102
rect 95294 274046 95362 274102
rect 95418 274046 125958 274102
rect 126014 274046 126082 274102
rect 126138 274046 156678 274102
rect 156734 274046 156802 274102
rect 156858 274046 187398 274102
rect 187454 274046 187522 274102
rect 187578 274046 218118 274102
rect 218174 274046 218242 274102
rect 218298 274046 248838 274102
rect 248894 274046 248962 274102
rect 249018 274046 279558 274102
rect 279614 274046 279682 274102
rect 279738 274046 310278 274102
rect 310334 274046 310402 274102
rect 310458 274046 340998 274102
rect 341054 274046 341122 274102
rect 341178 274046 363250 274102
rect 363306 274046 363374 274102
rect 363430 274046 363498 274102
rect 363554 274046 363622 274102
rect 363678 274046 371718 274102
rect 371774 274046 371842 274102
rect 371898 274046 381250 274102
rect 381306 274046 381374 274102
rect 381430 274046 381498 274102
rect 381554 274046 381622 274102
rect 381678 274046 399250 274102
rect 399306 274046 399374 274102
rect 399430 274046 399498 274102
rect 399554 274046 399622 274102
rect 399678 274046 402438 274102
rect 402494 274046 402562 274102
rect 402618 274046 433158 274102
rect 433214 274046 433282 274102
rect 433338 274046 435250 274102
rect 435306 274046 435374 274102
rect 435430 274046 435498 274102
rect 435554 274046 435622 274102
rect 435678 274046 453250 274102
rect 453306 274046 453374 274102
rect 453430 274046 453498 274102
rect 453554 274046 453622 274102
rect 453678 274046 471250 274102
rect 471306 274046 471374 274102
rect 471430 274046 471498 274102
rect 471554 274046 471622 274102
rect 471678 274046 489250 274102
rect 489306 274046 489374 274102
rect 489430 274046 489498 274102
rect 489554 274046 489622 274102
rect 489678 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 64518 273978
rect 64574 273922 64642 273978
rect 64698 273922 95238 273978
rect 95294 273922 95362 273978
rect 95418 273922 125958 273978
rect 126014 273922 126082 273978
rect 126138 273922 156678 273978
rect 156734 273922 156802 273978
rect 156858 273922 187398 273978
rect 187454 273922 187522 273978
rect 187578 273922 218118 273978
rect 218174 273922 218242 273978
rect 218298 273922 248838 273978
rect 248894 273922 248962 273978
rect 249018 273922 279558 273978
rect 279614 273922 279682 273978
rect 279738 273922 310278 273978
rect 310334 273922 310402 273978
rect 310458 273922 340998 273978
rect 341054 273922 341122 273978
rect 341178 273922 363250 273978
rect 363306 273922 363374 273978
rect 363430 273922 363498 273978
rect 363554 273922 363622 273978
rect 363678 273922 371718 273978
rect 371774 273922 371842 273978
rect 371898 273922 381250 273978
rect 381306 273922 381374 273978
rect 381430 273922 381498 273978
rect 381554 273922 381622 273978
rect 381678 273922 399250 273978
rect 399306 273922 399374 273978
rect 399430 273922 399498 273978
rect 399554 273922 399622 273978
rect 399678 273922 402438 273978
rect 402494 273922 402562 273978
rect 402618 273922 433158 273978
rect 433214 273922 433282 273978
rect 433338 273922 435250 273978
rect 435306 273922 435374 273978
rect 435430 273922 435498 273978
rect 435554 273922 435622 273978
rect 435678 273922 453250 273978
rect 453306 273922 453374 273978
rect 453430 273922 453498 273978
rect 453554 273922 453622 273978
rect 453678 273922 471250 273978
rect 471306 273922 471374 273978
rect 471430 273922 471498 273978
rect 471554 273922 471622 273978
rect 471678 273922 489250 273978
rect 489306 273922 489374 273978
rect 489430 273922 489498 273978
rect 489554 273922 489622 273978
rect 489678 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 79878 262350
rect 79934 262294 80002 262350
rect 80058 262294 110598 262350
rect 110654 262294 110722 262350
rect 110778 262294 141318 262350
rect 141374 262294 141442 262350
rect 141498 262294 172038 262350
rect 172094 262294 172162 262350
rect 172218 262294 202758 262350
rect 202814 262294 202882 262350
rect 202938 262294 233478 262350
rect 233534 262294 233602 262350
rect 233658 262294 264198 262350
rect 264254 262294 264322 262350
rect 264378 262294 294918 262350
rect 294974 262294 295042 262350
rect 295098 262294 325638 262350
rect 325694 262294 325762 262350
rect 325818 262294 348970 262350
rect 349026 262294 349094 262350
rect 349150 262294 349218 262350
rect 349274 262294 349342 262350
rect 349398 262294 356358 262350
rect 356414 262294 356482 262350
rect 356538 262294 366970 262350
rect 367026 262294 367094 262350
rect 367150 262294 367218 262350
rect 367274 262294 367342 262350
rect 367398 262294 384970 262350
rect 385026 262294 385094 262350
rect 385150 262294 385218 262350
rect 385274 262294 385342 262350
rect 385398 262294 387078 262350
rect 387134 262294 387202 262350
rect 387258 262294 402970 262350
rect 403026 262294 403094 262350
rect 403150 262294 403218 262350
rect 403274 262294 403342 262350
rect 403398 262294 417798 262350
rect 417854 262294 417922 262350
rect 417978 262294 420970 262350
rect 421026 262294 421094 262350
rect 421150 262294 421218 262350
rect 421274 262294 421342 262350
rect 421398 262294 438970 262350
rect 439026 262294 439094 262350
rect 439150 262294 439218 262350
rect 439274 262294 439342 262350
rect 439398 262294 456970 262350
rect 457026 262294 457094 262350
rect 457150 262294 457218 262350
rect 457274 262294 457342 262350
rect 457398 262294 474970 262350
rect 475026 262294 475094 262350
rect 475150 262294 475218 262350
rect 475274 262294 475342 262350
rect 475398 262294 492970 262350
rect 493026 262294 493094 262350
rect 493150 262294 493218 262350
rect 493274 262294 493342 262350
rect 493398 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 79878 262226
rect 79934 262170 80002 262226
rect 80058 262170 110598 262226
rect 110654 262170 110722 262226
rect 110778 262170 141318 262226
rect 141374 262170 141442 262226
rect 141498 262170 172038 262226
rect 172094 262170 172162 262226
rect 172218 262170 202758 262226
rect 202814 262170 202882 262226
rect 202938 262170 233478 262226
rect 233534 262170 233602 262226
rect 233658 262170 264198 262226
rect 264254 262170 264322 262226
rect 264378 262170 294918 262226
rect 294974 262170 295042 262226
rect 295098 262170 325638 262226
rect 325694 262170 325762 262226
rect 325818 262170 348970 262226
rect 349026 262170 349094 262226
rect 349150 262170 349218 262226
rect 349274 262170 349342 262226
rect 349398 262170 356358 262226
rect 356414 262170 356482 262226
rect 356538 262170 366970 262226
rect 367026 262170 367094 262226
rect 367150 262170 367218 262226
rect 367274 262170 367342 262226
rect 367398 262170 384970 262226
rect 385026 262170 385094 262226
rect 385150 262170 385218 262226
rect 385274 262170 385342 262226
rect 385398 262170 387078 262226
rect 387134 262170 387202 262226
rect 387258 262170 402970 262226
rect 403026 262170 403094 262226
rect 403150 262170 403218 262226
rect 403274 262170 403342 262226
rect 403398 262170 417798 262226
rect 417854 262170 417922 262226
rect 417978 262170 420970 262226
rect 421026 262170 421094 262226
rect 421150 262170 421218 262226
rect 421274 262170 421342 262226
rect 421398 262170 438970 262226
rect 439026 262170 439094 262226
rect 439150 262170 439218 262226
rect 439274 262170 439342 262226
rect 439398 262170 456970 262226
rect 457026 262170 457094 262226
rect 457150 262170 457218 262226
rect 457274 262170 457342 262226
rect 457398 262170 474970 262226
rect 475026 262170 475094 262226
rect 475150 262170 475218 262226
rect 475274 262170 475342 262226
rect 475398 262170 492970 262226
rect 493026 262170 493094 262226
rect 493150 262170 493218 262226
rect 493274 262170 493342 262226
rect 493398 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 79878 262102
rect 79934 262046 80002 262102
rect 80058 262046 110598 262102
rect 110654 262046 110722 262102
rect 110778 262046 141318 262102
rect 141374 262046 141442 262102
rect 141498 262046 172038 262102
rect 172094 262046 172162 262102
rect 172218 262046 202758 262102
rect 202814 262046 202882 262102
rect 202938 262046 233478 262102
rect 233534 262046 233602 262102
rect 233658 262046 264198 262102
rect 264254 262046 264322 262102
rect 264378 262046 294918 262102
rect 294974 262046 295042 262102
rect 295098 262046 325638 262102
rect 325694 262046 325762 262102
rect 325818 262046 348970 262102
rect 349026 262046 349094 262102
rect 349150 262046 349218 262102
rect 349274 262046 349342 262102
rect 349398 262046 356358 262102
rect 356414 262046 356482 262102
rect 356538 262046 366970 262102
rect 367026 262046 367094 262102
rect 367150 262046 367218 262102
rect 367274 262046 367342 262102
rect 367398 262046 384970 262102
rect 385026 262046 385094 262102
rect 385150 262046 385218 262102
rect 385274 262046 385342 262102
rect 385398 262046 387078 262102
rect 387134 262046 387202 262102
rect 387258 262046 402970 262102
rect 403026 262046 403094 262102
rect 403150 262046 403218 262102
rect 403274 262046 403342 262102
rect 403398 262046 417798 262102
rect 417854 262046 417922 262102
rect 417978 262046 420970 262102
rect 421026 262046 421094 262102
rect 421150 262046 421218 262102
rect 421274 262046 421342 262102
rect 421398 262046 438970 262102
rect 439026 262046 439094 262102
rect 439150 262046 439218 262102
rect 439274 262046 439342 262102
rect 439398 262046 456970 262102
rect 457026 262046 457094 262102
rect 457150 262046 457218 262102
rect 457274 262046 457342 262102
rect 457398 262046 474970 262102
rect 475026 262046 475094 262102
rect 475150 262046 475218 262102
rect 475274 262046 475342 262102
rect 475398 262046 492970 262102
rect 493026 262046 493094 262102
rect 493150 262046 493218 262102
rect 493274 262046 493342 262102
rect 493398 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 79878 261978
rect 79934 261922 80002 261978
rect 80058 261922 110598 261978
rect 110654 261922 110722 261978
rect 110778 261922 141318 261978
rect 141374 261922 141442 261978
rect 141498 261922 172038 261978
rect 172094 261922 172162 261978
rect 172218 261922 202758 261978
rect 202814 261922 202882 261978
rect 202938 261922 233478 261978
rect 233534 261922 233602 261978
rect 233658 261922 264198 261978
rect 264254 261922 264322 261978
rect 264378 261922 294918 261978
rect 294974 261922 295042 261978
rect 295098 261922 325638 261978
rect 325694 261922 325762 261978
rect 325818 261922 348970 261978
rect 349026 261922 349094 261978
rect 349150 261922 349218 261978
rect 349274 261922 349342 261978
rect 349398 261922 356358 261978
rect 356414 261922 356482 261978
rect 356538 261922 366970 261978
rect 367026 261922 367094 261978
rect 367150 261922 367218 261978
rect 367274 261922 367342 261978
rect 367398 261922 384970 261978
rect 385026 261922 385094 261978
rect 385150 261922 385218 261978
rect 385274 261922 385342 261978
rect 385398 261922 387078 261978
rect 387134 261922 387202 261978
rect 387258 261922 402970 261978
rect 403026 261922 403094 261978
rect 403150 261922 403218 261978
rect 403274 261922 403342 261978
rect 403398 261922 417798 261978
rect 417854 261922 417922 261978
rect 417978 261922 420970 261978
rect 421026 261922 421094 261978
rect 421150 261922 421218 261978
rect 421274 261922 421342 261978
rect 421398 261922 438970 261978
rect 439026 261922 439094 261978
rect 439150 261922 439218 261978
rect 439274 261922 439342 261978
rect 439398 261922 456970 261978
rect 457026 261922 457094 261978
rect 457150 261922 457218 261978
rect 457274 261922 457342 261978
rect 457398 261922 474970 261978
rect 475026 261922 475094 261978
rect 475150 261922 475218 261978
rect 475274 261922 475342 261978
rect 475398 261922 492970 261978
rect 493026 261922 493094 261978
rect 493150 261922 493218 261978
rect 493274 261922 493342 261978
rect 493398 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 64518 256350
rect 64574 256294 64642 256350
rect 64698 256294 95238 256350
rect 95294 256294 95362 256350
rect 95418 256294 125958 256350
rect 126014 256294 126082 256350
rect 126138 256294 156678 256350
rect 156734 256294 156802 256350
rect 156858 256294 187398 256350
rect 187454 256294 187522 256350
rect 187578 256294 218118 256350
rect 218174 256294 218242 256350
rect 218298 256294 248838 256350
rect 248894 256294 248962 256350
rect 249018 256294 279558 256350
rect 279614 256294 279682 256350
rect 279738 256294 310278 256350
rect 310334 256294 310402 256350
rect 310458 256294 340998 256350
rect 341054 256294 341122 256350
rect 341178 256294 363250 256350
rect 363306 256294 363374 256350
rect 363430 256294 363498 256350
rect 363554 256294 363622 256350
rect 363678 256294 371718 256350
rect 371774 256294 371842 256350
rect 371898 256294 381250 256350
rect 381306 256294 381374 256350
rect 381430 256294 381498 256350
rect 381554 256294 381622 256350
rect 381678 256294 399250 256350
rect 399306 256294 399374 256350
rect 399430 256294 399498 256350
rect 399554 256294 399622 256350
rect 399678 256294 402438 256350
rect 402494 256294 402562 256350
rect 402618 256294 433158 256350
rect 433214 256294 433282 256350
rect 433338 256294 435250 256350
rect 435306 256294 435374 256350
rect 435430 256294 435498 256350
rect 435554 256294 435622 256350
rect 435678 256294 453250 256350
rect 453306 256294 453374 256350
rect 453430 256294 453498 256350
rect 453554 256294 453622 256350
rect 453678 256294 471250 256350
rect 471306 256294 471374 256350
rect 471430 256294 471498 256350
rect 471554 256294 471622 256350
rect 471678 256294 489250 256350
rect 489306 256294 489374 256350
rect 489430 256294 489498 256350
rect 489554 256294 489622 256350
rect 489678 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 64518 256226
rect 64574 256170 64642 256226
rect 64698 256170 95238 256226
rect 95294 256170 95362 256226
rect 95418 256170 125958 256226
rect 126014 256170 126082 256226
rect 126138 256170 156678 256226
rect 156734 256170 156802 256226
rect 156858 256170 187398 256226
rect 187454 256170 187522 256226
rect 187578 256170 218118 256226
rect 218174 256170 218242 256226
rect 218298 256170 248838 256226
rect 248894 256170 248962 256226
rect 249018 256170 279558 256226
rect 279614 256170 279682 256226
rect 279738 256170 310278 256226
rect 310334 256170 310402 256226
rect 310458 256170 340998 256226
rect 341054 256170 341122 256226
rect 341178 256170 363250 256226
rect 363306 256170 363374 256226
rect 363430 256170 363498 256226
rect 363554 256170 363622 256226
rect 363678 256170 371718 256226
rect 371774 256170 371842 256226
rect 371898 256170 381250 256226
rect 381306 256170 381374 256226
rect 381430 256170 381498 256226
rect 381554 256170 381622 256226
rect 381678 256170 399250 256226
rect 399306 256170 399374 256226
rect 399430 256170 399498 256226
rect 399554 256170 399622 256226
rect 399678 256170 402438 256226
rect 402494 256170 402562 256226
rect 402618 256170 433158 256226
rect 433214 256170 433282 256226
rect 433338 256170 435250 256226
rect 435306 256170 435374 256226
rect 435430 256170 435498 256226
rect 435554 256170 435622 256226
rect 435678 256170 453250 256226
rect 453306 256170 453374 256226
rect 453430 256170 453498 256226
rect 453554 256170 453622 256226
rect 453678 256170 471250 256226
rect 471306 256170 471374 256226
rect 471430 256170 471498 256226
rect 471554 256170 471622 256226
rect 471678 256170 489250 256226
rect 489306 256170 489374 256226
rect 489430 256170 489498 256226
rect 489554 256170 489622 256226
rect 489678 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 64518 256102
rect 64574 256046 64642 256102
rect 64698 256046 95238 256102
rect 95294 256046 95362 256102
rect 95418 256046 125958 256102
rect 126014 256046 126082 256102
rect 126138 256046 156678 256102
rect 156734 256046 156802 256102
rect 156858 256046 187398 256102
rect 187454 256046 187522 256102
rect 187578 256046 218118 256102
rect 218174 256046 218242 256102
rect 218298 256046 248838 256102
rect 248894 256046 248962 256102
rect 249018 256046 279558 256102
rect 279614 256046 279682 256102
rect 279738 256046 310278 256102
rect 310334 256046 310402 256102
rect 310458 256046 340998 256102
rect 341054 256046 341122 256102
rect 341178 256046 363250 256102
rect 363306 256046 363374 256102
rect 363430 256046 363498 256102
rect 363554 256046 363622 256102
rect 363678 256046 371718 256102
rect 371774 256046 371842 256102
rect 371898 256046 381250 256102
rect 381306 256046 381374 256102
rect 381430 256046 381498 256102
rect 381554 256046 381622 256102
rect 381678 256046 399250 256102
rect 399306 256046 399374 256102
rect 399430 256046 399498 256102
rect 399554 256046 399622 256102
rect 399678 256046 402438 256102
rect 402494 256046 402562 256102
rect 402618 256046 433158 256102
rect 433214 256046 433282 256102
rect 433338 256046 435250 256102
rect 435306 256046 435374 256102
rect 435430 256046 435498 256102
rect 435554 256046 435622 256102
rect 435678 256046 453250 256102
rect 453306 256046 453374 256102
rect 453430 256046 453498 256102
rect 453554 256046 453622 256102
rect 453678 256046 471250 256102
rect 471306 256046 471374 256102
rect 471430 256046 471498 256102
rect 471554 256046 471622 256102
rect 471678 256046 489250 256102
rect 489306 256046 489374 256102
rect 489430 256046 489498 256102
rect 489554 256046 489622 256102
rect 489678 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 64518 255978
rect 64574 255922 64642 255978
rect 64698 255922 95238 255978
rect 95294 255922 95362 255978
rect 95418 255922 125958 255978
rect 126014 255922 126082 255978
rect 126138 255922 156678 255978
rect 156734 255922 156802 255978
rect 156858 255922 187398 255978
rect 187454 255922 187522 255978
rect 187578 255922 218118 255978
rect 218174 255922 218242 255978
rect 218298 255922 248838 255978
rect 248894 255922 248962 255978
rect 249018 255922 279558 255978
rect 279614 255922 279682 255978
rect 279738 255922 310278 255978
rect 310334 255922 310402 255978
rect 310458 255922 340998 255978
rect 341054 255922 341122 255978
rect 341178 255922 363250 255978
rect 363306 255922 363374 255978
rect 363430 255922 363498 255978
rect 363554 255922 363622 255978
rect 363678 255922 371718 255978
rect 371774 255922 371842 255978
rect 371898 255922 381250 255978
rect 381306 255922 381374 255978
rect 381430 255922 381498 255978
rect 381554 255922 381622 255978
rect 381678 255922 399250 255978
rect 399306 255922 399374 255978
rect 399430 255922 399498 255978
rect 399554 255922 399622 255978
rect 399678 255922 402438 255978
rect 402494 255922 402562 255978
rect 402618 255922 433158 255978
rect 433214 255922 433282 255978
rect 433338 255922 435250 255978
rect 435306 255922 435374 255978
rect 435430 255922 435498 255978
rect 435554 255922 435622 255978
rect 435678 255922 453250 255978
rect 453306 255922 453374 255978
rect 453430 255922 453498 255978
rect 453554 255922 453622 255978
rect 453678 255922 471250 255978
rect 471306 255922 471374 255978
rect 471430 255922 471498 255978
rect 471554 255922 471622 255978
rect 471678 255922 489250 255978
rect 489306 255922 489374 255978
rect 489430 255922 489498 255978
rect 489554 255922 489622 255978
rect 489678 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 79878 244350
rect 79934 244294 80002 244350
rect 80058 244294 110598 244350
rect 110654 244294 110722 244350
rect 110778 244294 141318 244350
rect 141374 244294 141442 244350
rect 141498 244294 172038 244350
rect 172094 244294 172162 244350
rect 172218 244294 202758 244350
rect 202814 244294 202882 244350
rect 202938 244294 233478 244350
rect 233534 244294 233602 244350
rect 233658 244294 264198 244350
rect 264254 244294 264322 244350
rect 264378 244294 294918 244350
rect 294974 244294 295042 244350
rect 295098 244294 325638 244350
rect 325694 244294 325762 244350
rect 325818 244294 348970 244350
rect 349026 244294 349094 244350
rect 349150 244294 349218 244350
rect 349274 244294 349342 244350
rect 349398 244294 356358 244350
rect 356414 244294 356482 244350
rect 356538 244294 366970 244350
rect 367026 244294 367094 244350
rect 367150 244294 367218 244350
rect 367274 244294 367342 244350
rect 367398 244294 384970 244350
rect 385026 244294 385094 244350
rect 385150 244294 385218 244350
rect 385274 244294 385342 244350
rect 385398 244294 387078 244350
rect 387134 244294 387202 244350
rect 387258 244294 402970 244350
rect 403026 244294 403094 244350
rect 403150 244294 403218 244350
rect 403274 244294 403342 244350
rect 403398 244294 417798 244350
rect 417854 244294 417922 244350
rect 417978 244294 420970 244350
rect 421026 244294 421094 244350
rect 421150 244294 421218 244350
rect 421274 244294 421342 244350
rect 421398 244294 438970 244350
rect 439026 244294 439094 244350
rect 439150 244294 439218 244350
rect 439274 244294 439342 244350
rect 439398 244294 456970 244350
rect 457026 244294 457094 244350
rect 457150 244294 457218 244350
rect 457274 244294 457342 244350
rect 457398 244294 474970 244350
rect 475026 244294 475094 244350
rect 475150 244294 475218 244350
rect 475274 244294 475342 244350
rect 475398 244294 492970 244350
rect 493026 244294 493094 244350
rect 493150 244294 493218 244350
rect 493274 244294 493342 244350
rect 493398 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 79878 244226
rect 79934 244170 80002 244226
rect 80058 244170 110598 244226
rect 110654 244170 110722 244226
rect 110778 244170 141318 244226
rect 141374 244170 141442 244226
rect 141498 244170 172038 244226
rect 172094 244170 172162 244226
rect 172218 244170 202758 244226
rect 202814 244170 202882 244226
rect 202938 244170 233478 244226
rect 233534 244170 233602 244226
rect 233658 244170 264198 244226
rect 264254 244170 264322 244226
rect 264378 244170 294918 244226
rect 294974 244170 295042 244226
rect 295098 244170 325638 244226
rect 325694 244170 325762 244226
rect 325818 244170 348970 244226
rect 349026 244170 349094 244226
rect 349150 244170 349218 244226
rect 349274 244170 349342 244226
rect 349398 244170 356358 244226
rect 356414 244170 356482 244226
rect 356538 244170 366970 244226
rect 367026 244170 367094 244226
rect 367150 244170 367218 244226
rect 367274 244170 367342 244226
rect 367398 244170 384970 244226
rect 385026 244170 385094 244226
rect 385150 244170 385218 244226
rect 385274 244170 385342 244226
rect 385398 244170 387078 244226
rect 387134 244170 387202 244226
rect 387258 244170 402970 244226
rect 403026 244170 403094 244226
rect 403150 244170 403218 244226
rect 403274 244170 403342 244226
rect 403398 244170 417798 244226
rect 417854 244170 417922 244226
rect 417978 244170 420970 244226
rect 421026 244170 421094 244226
rect 421150 244170 421218 244226
rect 421274 244170 421342 244226
rect 421398 244170 438970 244226
rect 439026 244170 439094 244226
rect 439150 244170 439218 244226
rect 439274 244170 439342 244226
rect 439398 244170 456970 244226
rect 457026 244170 457094 244226
rect 457150 244170 457218 244226
rect 457274 244170 457342 244226
rect 457398 244170 474970 244226
rect 475026 244170 475094 244226
rect 475150 244170 475218 244226
rect 475274 244170 475342 244226
rect 475398 244170 492970 244226
rect 493026 244170 493094 244226
rect 493150 244170 493218 244226
rect 493274 244170 493342 244226
rect 493398 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 79878 244102
rect 79934 244046 80002 244102
rect 80058 244046 110598 244102
rect 110654 244046 110722 244102
rect 110778 244046 141318 244102
rect 141374 244046 141442 244102
rect 141498 244046 172038 244102
rect 172094 244046 172162 244102
rect 172218 244046 202758 244102
rect 202814 244046 202882 244102
rect 202938 244046 233478 244102
rect 233534 244046 233602 244102
rect 233658 244046 264198 244102
rect 264254 244046 264322 244102
rect 264378 244046 294918 244102
rect 294974 244046 295042 244102
rect 295098 244046 325638 244102
rect 325694 244046 325762 244102
rect 325818 244046 348970 244102
rect 349026 244046 349094 244102
rect 349150 244046 349218 244102
rect 349274 244046 349342 244102
rect 349398 244046 356358 244102
rect 356414 244046 356482 244102
rect 356538 244046 366970 244102
rect 367026 244046 367094 244102
rect 367150 244046 367218 244102
rect 367274 244046 367342 244102
rect 367398 244046 384970 244102
rect 385026 244046 385094 244102
rect 385150 244046 385218 244102
rect 385274 244046 385342 244102
rect 385398 244046 387078 244102
rect 387134 244046 387202 244102
rect 387258 244046 402970 244102
rect 403026 244046 403094 244102
rect 403150 244046 403218 244102
rect 403274 244046 403342 244102
rect 403398 244046 417798 244102
rect 417854 244046 417922 244102
rect 417978 244046 420970 244102
rect 421026 244046 421094 244102
rect 421150 244046 421218 244102
rect 421274 244046 421342 244102
rect 421398 244046 438970 244102
rect 439026 244046 439094 244102
rect 439150 244046 439218 244102
rect 439274 244046 439342 244102
rect 439398 244046 456970 244102
rect 457026 244046 457094 244102
rect 457150 244046 457218 244102
rect 457274 244046 457342 244102
rect 457398 244046 474970 244102
rect 475026 244046 475094 244102
rect 475150 244046 475218 244102
rect 475274 244046 475342 244102
rect 475398 244046 492970 244102
rect 493026 244046 493094 244102
rect 493150 244046 493218 244102
rect 493274 244046 493342 244102
rect 493398 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 79878 243978
rect 79934 243922 80002 243978
rect 80058 243922 110598 243978
rect 110654 243922 110722 243978
rect 110778 243922 141318 243978
rect 141374 243922 141442 243978
rect 141498 243922 172038 243978
rect 172094 243922 172162 243978
rect 172218 243922 202758 243978
rect 202814 243922 202882 243978
rect 202938 243922 233478 243978
rect 233534 243922 233602 243978
rect 233658 243922 264198 243978
rect 264254 243922 264322 243978
rect 264378 243922 294918 243978
rect 294974 243922 295042 243978
rect 295098 243922 325638 243978
rect 325694 243922 325762 243978
rect 325818 243922 348970 243978
rect 349026 243922 349094 243978
rect 349150 243922 349218 243978
rect 349274 243922 349342 243978
rect 349398 243922 356358 243978
rect 356414 243922 356482 243978
rect 356538 243922 366970 243978
rect 367026 243922 367094 243978
rect 367150 243922 367218 243978
rect 367274 243922 367342 243978
rect 367398 243922 384970 243978
rect 385026 243922 385094 243978
rect 385150 243922 385218 243978
rect 385274 243922 385342 243978
rect 385398 243922 387078 243978
rect 387134 243922 387202 243978
rect 387258 243922 402970 243978
rect 403026 243922 403094 243978
rect 403150 243922 403218 243978
rect 403274 243922 403342 243978
rect 403398 243922 417798 243978
rect 417854 243922 417922 243978
rect 417978 243922 420970 243978
rect 421026 243922 421094 243978
rect 421150 243922 421218 243978
rect 421274 243922 421342 243978
rect 421398 243922 438970 243978
rect 439026 243922 439094 243978
rect 439150 243922 439218 243978
rect 439274 243922 439342 243978
rect 439398 243922 456970 243978
rect 457026 243922 457094 243978
rect 457150 243922 457218 243978
rect 457274 243922 457342 243978
rect 457398 243922 474970 243978
rect 475026 243922 475094 243978
rect 475150 243922 475218 243978
rect 475274 243922 475342 243978
rect 475398 243922 492970 243978
rect 493026 243922 493094 243978
rect 493150 243922 493218 243978
rect 493274 243922 493342 243978
rect 493398 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 64518 238350
rect 64574 238294 64642 238350
rect 64698 238294 95238 238350
rect 95294 238294 95362 238350
rect 95418 238294 125958 238350
rect 126014 238294 126082 238350
rect 126138 238294 156678 238350
rect 156734 238294 156802 238350
rect 156858 238294 187398 238350
rect 187454 238294 187522 238350
rect 187578 238294 218118 238350
rect 218174 238294 218242 238350
rect 218298 238294 248838 238350
rect 248894 238294 248962 238350
rect 249018 238294 279558 238350
rect 279614 238294 279682 238350
rect 279738 238294 310278 238350
rect 310334 238294 310402 238350
rect 310458 238294 340998 238350
rect 341054 238294 341122 238350
rect 341178 238294 363250 238350
rect 363306 238294 363374 238350
rect 363430 238294 363498 238350
rect 363554 238294 363622 238350
rect 363678 238294 371718 238350
rect 371774 238294 371842 238350
rect 371898 238294 381250 238350
rect 381306 238294 381374 238350
rect 381430 238294 381498 238350
rect 381554 238294 381622 238350
rect 381678 238294 399250 238350
rect 399306 238294 399374 238350
rect 399430 238294 399498 238350
rect 399554 238294 399622 238350
rect 399678 238294 402438 238350
rect 402494 238294 402562 238350
rect 402618 238294 433158 238350
rect 433214 238294 433282 238350
rect 433338 238294 435250 238350
rect 435306 238294 435374 238350
rect 435430 238294 435498 238350
rect 435554 238294 435622 238350
rect 435678 238294 453250 238350
rect 453306 238294 453374 238350
rect 453430 238294 453498 238350
rect 453554 238294 453622 238350
rect 453678 238294 471250 238350
rect 471306 238294 471374 238350
rect 471430 238294 471498 238350
rect 471554 238294 471622 238350
rect 471678 238294 489250 238350
rect 489306 238294 489374 238350
rect 489430 238294 489498 238350
rect 489554 238294 489622 238350
rect 489678 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 64518 238226
rect 64574 238170 64642 238226
rect 64698 238170 95238 238226
rect 95294 238170 95362 238226
rect 95418 238170 125958 238226
rect 126014 238170 126082 238226
rect 126138 238170 156678 238226
rect 156734 238170 156802 238226
rect 156858 238170 187398 238226
rect 187454 238170 187522 238226
rect 187578 238170 218118 238226
rect 218174 238170 218242 238226
rect 218298 238170 248838 238226
rect 248894 238170 248962 238226
rect 249018 238170 279558 238226
rect 279614 238170 279682 238226
rect 279738 238170 310278 238226
rect 310334 238170 310402 238226
rect 310458 238170 340998 238226
rect 341054 238170 341122 238226
rect 341178 238170 363250 238226
rect 363306 238170 363374 238226
rect 363430 238170 363498 238226
rect 363554 238170 363622 238226
rect 363678 238170 371718 238226
rect 371774 238170 371842 238226
rect 371898 238170 381250 238226
rect 381306 238170 381374 238226
rect 381430 238170 381498 238226
rect 381554 238170 381622 238226
rect 381678 238170 399250 238226
rect 399306 238170 399374 238226
rect 399430 238170 399498 238226
rect 399554 238170 399622 238226
rect 399678 238170 402438 238226
rect 402494 238170 402562 238226
rect 402618 238170 433158 238226
rect 433214 238170 433282 238226
rect 433338 238170 435250 238226
rect 435306 238170 435374 238226
rect 435430 238170 435498 238226
rect 435554 238170 435622 238226
rect 435678 238170 453250 238226
rect 453306 238170 453374 238226
rect 453430 238170 453498 238226
rect 453554 238170 453622 238226
rect 453678 238170 471250 238226
rect 471306 238170 471374 238226
rect 471430 238170 471498 238226
rect 471554 238170 471622 238226
rect 471678 238170 489250 238226
rect 489306 238170 489374 238226
rect 489430 238170 489498 238226
rect 489554 238170 489622 238226
rect 489678 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 64518 238102
rect 64574 238046 64642 238102
rect 64698 238046 95238 238102
rect 95294 238046 95362 238102
rect 95418 238046 125958 238102
rect 126014 238046 126082 238102
rect 126138 238046 156678 238102
rect 156734 238046 156802 238102
rect 156858 238046 187398 238102
rect 187454 238046 187522 238102
rect 187578 238046 218118 238102
rect 218174 238046 218242 238102
rect 218298 238046 248838 238102
rect 248894 238046 248962 238102
rect 249018 238046 279558 238102
rect 279614 238046 279682 238102
rect 279738 238046 310278 238102
rect 310334 238046 310402 238102
rect 310458 238046 340998 238102
rect 341054 238046 341122 238102
rect 341178 238046 363250 238102
rect 363306 238046 363374 238102
rect 363430 238046 363498 238102
rect 363554 238046 363622 238102
rect 363678 238046 371718 238102
rect 371774 238046 371842 238102
rect 371898 238046 381250 238102
rect 381306 238046 381374 238102
rect 381430 238046 381498 238102
rect 381554 238046 381622 238102
rect 381678 238046 399250 238102
rect 399306 238046 399374 238102
rect 399430 238046 399498 238102
rect 399554 238046 399622 238102
rect 399678 238046 402438 238102
rect 402494 238046 402562 238102
rect 402618 238046 433158 238102
rect 433214 238046 433282 238102
rect 433338 238046 435250 238102
rect 435306 238046 435374 238102
rect 435430 238046 435498 238102
rect 435554 238046 435622 238102
rect 435678 238046 453250 238102
rect 453306 238046 453374 238102
rect 453430 238046 453498 238102
rect 453554 238046 453622 238102
rect 453678 238046 471250 238102
rect 471306 238046 471374 238102
rect 471430 238046 471498 238102
rect 471554 238046 471622 238102
rect 471678 238046 489250 238102
rect 489306 238046 489374 238102
rect 489430 238046 489498 238102
rect 489554 238046 489622 238102
rect 489678 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 64518 237978
rect 64574 237922 64642 237978
rect 64698 237922 95238 237978
rect 95294 237922 95362 237978
rect 95418 237922 125958 237978
rect 126014 237922 126082 237978
rect 126138 237922 156678 237978
rect 156734 237922 156802 237978
rect 156858 237922 187398 237978
rect 187454 237922 187522 237978
rect 187578 237922 218118 237978
rect 218174 237922 218242 237978
rect 218298 237922 248838 237978
rect 248894 237922 248962 237978
rect 249018 237922 279558 237978
rect 279614 237922 279682 237978
rect 279738 237922 310278 237978
rect 310334 237922 310402 237978
rect 310458 237922 340998 237978
rect 341054 237922 341122 237978
rect 341178 237922 363250 237978
rect 363306 237922 363374 237978
rect 363430 237922 363498 237978
rect 363554 237922 363622 237978
rect 363678 237922 371718 237978
rect 371774 237922 371842 237978
rect 371898 237922 381250 237978
rect 381306 237922 381374 237978
rect 381430 237922 381498 237978
rect 381554 237922 381622 237978
rect 381678 237922 399250 237978
rect 399306 237922 399374 237978
rect 399430 237922 399498 237978
rect 399554 237922 399622 237978
rect 399678 237922 402438 237978
rect 402494 237922 402562 237978
rect 402618 237922 433158 237978
rect 433214 237922 433282 237978
rect 433338 237922 435250 237978
rect 435306 237922 435374 237978
rect 435430 237922 435498 237978
rect 435554 237922 435622 237978
rect 435678 237922 453250 237978
rect 453306 237922 453374 237978
rect 453430 237922 453498 237978
rect 453554 237922 453622 237978
rect 453678 237922 471250 237978
rect 471306 237922 471374 237978
rect 471430 237922 471498 237978
rect 471554 237922 471622 237978
rect 471678 237922 489250 237978
rect 489306 237922 489374 237978
rect 489430 237922 489498 237978
rect 489554 237922 489622 237978
rect 489678 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 79878 226350
rect 79934 226294 80002 226350
rect 80058 226294 110598 226350
rect 110654 226294 110722 226350
rect 110778 226294 141318 226350
rect 141374 226294 141442 226350
rect 141498 226294 172038 226350
rect 172094 226294 172162 226350
rect 172218 226294 202758 226350
rect 202814 226294 202882 226350
rect 202938 226294 233478 226350
rect 233534 226294 233602 226350
rect 233658 226294 264198 226350
rect 264254 226294 264322 226350
rect 264378 226294 294918 226350
rect 294974 226294 295042 226350
rect 295098 226294 325638 226350
rect 325694 226294 325762 226350
rect 325818 226294 348970 226350
rect 349026 226294 349094 226350
rect 349150 226294 349218 226350
rect 349274 226294 349342 226350
rect 349398 226294 356358 226350
rect 356414 226294 356482 226350
rect 356538 226294 366970 226350
rect 367026 226294 367094 226350
rect 367150 226294 367218 226350
rect 367274 226294 367342 226350
rect 367398 226294 384970 226350
rect 385026 226294 385094 226350
rect 385150 226294 385218 226350
rect 385274 226294 385342 226350
rect 385398 226294 387078 226350
rect 387134 226294 387202 226350
rect 387258 226294 402970 226350
rect 403026 226294 403094 226350
rect 403150 226294 403218 226350
rect 403274 226294 403342 226350
rect 403398 226294 417798 226350
rect 417854 226294 417922 226350
rect 417978 226294 420970 226350
rect 421026 226294 421094 226350
rect 421150 226294 421218 226350
rect 421274 226294 421342 226350
rect 421398 226294 438970 226350
rect 439026 226294 439094 226350
rect 439150 226294 439218 226350
rect 439274 226294 439342 226350
rect 439398 226294 456970 226350
rect 457026 226294 457094 226350
rect 457150 226294 457218 226350
rect 457274 226294 457342 226350
rect 457398 226294 474970 226350
rect 475026 226294 475094 226350
rect 475150 226294 475218 226350
rect 475274 226294 475342 226350
rect 475398 226294 492970 226350
rect 493026 226294 493094 226350
rect 493150 226294 493218 226350
rect 493274 226294 493342 226350
rect 493398 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 79878 226226
rect 79934 226170 80002 226226
rect 80058 226170 110598 226226
rect 110654 226170 110722 226226
rect 110778 226170 141318 226226
rect 141374 226170 141442 226226
rect 141498 226170 172038 226226
rect 172094 226170 172162 226226
rect 172218 226170 202758 226226
rect 202814 226170 202882 226226
rect 202938 226170 233478 226226
rect 233534 226170 233602 226226
rect 233658 226170 264198 226226
rect 264254 226170 264322 226226
rect 264378 226170 294918 226226
rect 294974 226170 295042 226226
rect 295098 226170 325638 226226
rect 325694 226170 325762 226226
rect 325818 226170 348970 226226
rect 349026 226170 349094 226226
rect 349150 226170 349218 226226
rect 349274 226170 349342 226226
rect 349398 226170 356358 226226
rect 356414 226170 356482 226226
rect 356538 226170 366970 226226
rect 367026 226170 367094 226226
rect 367150 226170 367218 226226
rect 367274 226170 367342 226226
rect 367398 226170 384970 226226
rect 385026 226170 385094 226226
rect 385150 226170 385218 226226
rect 385274 226170 385342 226226
rect 385398 226170 387078 226226
rect 387134 226170 387202 226226
rect 387258 226170 402970 226226
rect 403026 226170 403094 226226
rect 403150 226170 403218 226226
rect 403274 226170 403342 226226
rect 403398 226170 417798 226226
rect 417854 226170 417922 226226
rect 417978 226170 420970 226226
rect 421026 226170 421094 226226
rect 421150 226170 421218 226226
rect 421274 226170 421342 226226
rect 421398 226170 438970 226226
rect 439026 226170 439094 226226
rect 439150 226170 439218 226226
rect 439274 226170 439342 226226
rect 439398 226170 456970 226226
rect 457026 226170 457094 226226
rect 457150 226170 457218 226226
rect 457274 226170 457342 226226
rect 457398 226170 474970 226226
rect 475026 226170 475094 226226
rect 475150 226170 475218 226226
rect 475274 226170 475342 226226
rect 475398 226170 492970 226226
rect 493026 226170 493094 226226
rect 493150 226170 493218 226226
rect 493274 226170 493342 226226
rect 493398 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 79878 226102
rect 79934 226046 80002 226102
rect 80058 226046 110598 226102
rect 110654 226046 110722 226102
rect 110778 226046 141318 226102
rect 141374 226046 141442 226102
rect 141498 226046 172038 226102
rect 172094 226046 172162 226102
rect 172218 226046 202758 226102
rect 202814 226046 202882 226102
rect 202938 226046 233478 226102
rect 233534 226046 233602 226102
rect 233658 226046 264198 226102
rect 264254 226046 264322 226102
rect 264378 226046 294918 226102
rect 294974 226046 295042 226102
rect 295098 226046 325638 226102
rect 325694 226046 325762 226102
rect 325818 226046 348970 226102
rect 349026 226046 349094 226102
rect 349150 226046 349218 226102
rect 349274 226046 349342 226102
rect 349398 226046 356358 226102
rect 356414 226046 356482 226102
rect 356538 226046 366970 226102
rect 367026 226046 367094 226102
rect 367150 226046 367218 226102
rect 367274 226046 367342 226102
rect 367398 226046 384970 226102
rect 385026 226046 385094 226102
rect 385150 226046 385218 226102
rect 385274 226046 385342 226102
rect 385398 226046 387078 226102
rect 387134 226046 387202 226102
rect 387258 226046 402970 226102
rect 403026 226046 403094 226102
rect 403150 226046 403218 226102
rect 403274 226046 403342 226102
rect 403398 226046 417798 226102
rect 417854 226046 417922 226102
rect 417978 226046 420970 226102
rect 421026 226046 421094 226102
rect 421150 226046 421218 226102
rect 421274 226046 421342 226102
rect 421398 226046 438970 226102
rect 439026 226046 439094 226102
rect 439150 226046 439218 226102
rect 439274 226046 439342 226102
rect 439398 226046 456970 226102
rect 457026 226046 457094 226102
rect 457150 226046 457218 226102
rect 457274 226046 457342 226102
rect 457398 226046 474970 226102
rect 475026 226046 475094 226102
rect 475150 226046 475218 226102
rect 475274 226046 475342 226102
rect 475398 226046 492970 226102
rect 493026 226046 493094 226102
rect 493150 226046 493218 226102
rect 493274 226046 493342 226102
rect 493398 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 79878 225978
rect 79934 225922 80002 225978
rect 80058 225922 110598 225978
rect 110654 225922 110722 225978
rect 110778 225922 141318 225978
rect 141374 225922 141442 225978
rect 141498 225922 172038 225978
rect 172094 225922 172162 225978
rect 172218 225922 202758 225978
rect 202814 225922 202882 225978
rect 202938 225922 233478 225978
rect 233534 225922 233602 225978
rect 233658 225922 264198 225978
rect 264254 225922 264322 225978
rect 264378 225922 294918 225978
rect 294974 225922 295042 225978
rect 295098 225922 325638 225978
rect 325694 225922 325762 225978
rect 325818 225922 348970 225978
rect 349026 225922 349094 225978
rect 349150 225922 349218 225978
rect 349274 225922 349342 225978
rect 349398 225922 356358 225978
rect 356414 225922 356482 225978
rect 356538 225922 366970 225978
rect 367026 225922 367094 225978
rect 367150 225922 367218 225978
rect 367274 225922 367342 225978
rect 367398 225922 384970 225978
rect 385026 225922 385094 225978
rect 385150 225922 385218 225978
rect 385274 225922 385342 225978
rect 385398 225922 387078 225978
rect 387134 225922 387202 225978
rect 387258 225922 402970 225978
rect 403026 225922 403094 225978
rect 403150 225922 403218 225978
rect 403274 225922 403342 225978
rect 403398 225922 417798 225978
rect 417854 225922 417922 225978
rect 417978 225922 420970 225978
rect 421026 225922 421094 225978
rect 421150 225922 421218 225978
rect 421274 225922 421342 225978
rect 421398 225922 438970 225978
rect 439026 225922 439094 225978
rect 439150 225922 439218 225978
rect 439274 225922 439342 225978
rect 439398 225922 456970 225978
rect 457026 225922 457094 225978
rect 457150 225922 457218 225978
rect 457274 225922 457342 225978
rect 457398 225922 474970 225978
rect 475026 225922 475094 225978
rect 475150 225922 475218 225978
rect 475274 225922 475342 225978
rect 475398 225922 492970 225978
rect 493026 225922 493094 225978
rect 493150 225922 493218 225978
rect 493274 225922 493342 225978
rect 493398 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 64518 220350
rect 64574 220294 64642 220350
rect 64698 220294 95238 220350
rect 95294 220294 95362 220350
rect 95418 220294 125958 220350
rect 126014 220294 126082 220350
rect 126138 220294 156678 220350
rect 156734 220294 156802 220350
rect 156858 220294 187398 220350
rect 187454 220294 187522 220350
rect 187578 220294 218118 220350
rect 218174 220294 218242 220350
rect 218298 220294 248838 220350
rect 248894 220294 248962 220350
rect 249018 220294 279558 220350
rect 279614 220294 279682 220350
rect 279738 220294 310278 220350
rect 310334 220294 310402 220350
rect 310458 220294 340998 220350
rect 341054 220294 341122 220350
rect 341178 220294 363250 220350
rect 363306 220294 363374 220350
rect 363430 220294 363498 220350
rect 363554 220294 363622 220350
rect 363678 220294 371718 220350
rect 371774 220294 371842 220350
rect 371898 220294 381250 220350
rect 381306 220294 381374 220350
rect 381430 220294 381498 220350
rect 381554 220294 381622 220350
rect 381678 220294 399250 220350
rect 399306 220294 399374 220350
rect 399430 220294 399498 220350
rect 399554 220294 399622 220350
rect 399678 220294 402438 220350
rect 402494 220294 402562 220350
rect 402618 220294 433158 220350
rect 433214 220294 433282 220350
rect 433338 220294 435250 220350
rect 435306 220294 435374 220350
rect 435430 220294 435498 220350
rect 435554 220294 435622 220350
rect 435678 220294 453250 220350
rect 453306 220294 453374 220350
rect 453430 220294 453498 220350
rect 453554 220294 453622 220350
rect 453678 220294 471250 220350
rect 471306 220294 471374 220350
rect 471430 220294 471498 220350
rect 471554 220294 471622 220350
rect 471678 220294 489250 220350
rect 489306 220294 489374 220350
rect 489430 220294 489498 220350
rect 489554 220294 489622 220350
rect 489678 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 64518 220226
rect 64574 220170 64642 220226
rect 64698 220170 95238 220226
rect 95294 220170 95362 220226
rect 95418 220170 125958 220226
rect 126014 220170 126082 220226
rect 126138 220170 156678 220226
rect 156734 220170 156802 220226
rect 156858 220170 187398 220226
rect 187454 220170 187522 220226
rect 187578 220170 218118 220226
rect 218174 220170 218242 220226
rect 218298 220170 248838 220226
rect 248894 220170 248962 220226
rect 249018 220170 279558 220226
rect 279614 220170 279682 220226
rect 279738 220170 310278 220226
rect 310334 220170 310402 220226
rect 310458 220170 340998 220226
rect 341054 220170 341122 220226
rect 341178 220170 363250 220226
rect 363306 220170 363374 220226
rect 363430 220170 363498 220226
rect 363554 220170 363622 220226
rect 363678 220170 371718 220226
rect 371774 220170 371842 220226
rect 371898 220170 381250 220226
rect 381306 220170 381374 220226
rect 381430 220170 381498 220226
rect 381554 220170 381622 220226
rect 381678 220170 399250 220226
rect 399306 220170 399374 220226
rect 399430 220170 399498 220226
rect 399554 220170 399622 220226
rect 399678 220170 402438 220226
rect 402494 220170 402562 220226
rect 402618 220170 433158 220226
rect 433214 220170 433282 220226
rect 433338 220170 435250 220226
rect 435306 220170 435374 220226
rect 435430 220170 435498 220226
rect 435554 220170 435622 220226
rect 435678 220170 453250 220226
rect 453306 220170 453374 220226
rect 453430 220170 453498 220226
rect 453554 220170 453622 220226
rect 453678 220170 471250 220226
rect 471306 220170 471374 220226
rect 471430 220170 471498 220226
rect 471554 220170 471622 220226
rect 471678 220170 489250 220226
rect 489306 220170 489374 220226
rect 489430 220170 489498 220226
rect 489554 220170 489622 220226
rect 489678 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 64518 220102
rect 64574 220046 64642 220102
rect 64698 220046 95238 220102
rect 95294 220046 95362 220102
rect 95418 220046 125958 220102
rect 126014 220046 126082 220102
rect 126138 220046 156678 220102
rect 156734 220046 156802 220102
rect 156858 220046 187398 220102
rect 187454 220046 187522 220102
rect 187578 220046 218118 220102
rect 218174 220046 218242 220102
rect 218298 220046 248838 220102
rect 248894 220046 248962 220102
rect 249018 220046 279558 220102
rect 279614 220046 279682 220102
rect 279738 220046 310278 220102
rect 310334 220046 310402 220102
rect 310458 220046 340998 220102
rect 341054 220046 341122 220102
rect 341178 220046 363250 220102
rect 363306 220046 363374 220102
rect 363430 220046 363498 220102
rect 363554 220046 363622 220102
rect 363678 220046 371718 220102
rect 371774 220046 371842 220102
rect 371898 220046 381250 220102
rect 381306 220046 381374 220102
rect 381430 220046 381498 220102
rect 381554 220046 381622 220102
rect 381678 220046 399250 220102
rect 399306 220046 399374 220102
rect 399430 220046 399498 220102
rect 399554 220046 399622 220102
rect 399678 220046 402438 220102
rect 402494 220046 402562 220102
rect 402618 220046 433158 220102
rect 433214 220046 433282 220102
rect 433338 220046 435250 220102
rect 435306 220046 435374 220102
rect 435430 220046 435498 220102
rect 435554 220046 435622 220102
rect 435678 220046 453250 220102
rect 453306 220046 453374 220102
rect 453430 220046 453498 220102
rect 453554 220046 453622 220102
rect 453678 220046 471250 220102
rect 471306 220046 471374 220102
rect 471430 220046 471498 220102
rect 471554 220046 471622 220102
rect 471678 220046 489250 220102
rect 489306 220046 489374 220102
rect 489430 220046 489498 220102
rect 489554 220046 489622 220102
rect 489678 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 64518 219978
rect 64574 219922 64642 219978
rect 64698 219922 95238 219978
rect 95294 219922 95362 219978
rect 95418 219922 125958 219978
rect 126014 219922 126082 219978
rect 126138 219922 156678 219978
rect 156734 219922 156802 219978
rect 156858 219922 187398 219978
rect 187454 219922 187522 219978
rect 187578 219922 218118 219978
rect 218174 219922 218242 219978
rect 218298 219922 248838 219978
rect 248894 219922 248962 219978
rect 249018 219922 279558 219978
rect 279614 219922 279682 219978
rect 279738 219922 310278 219978
rect 310334 219922 310402 219978
rect 310458 219922 340998 219978
rect 341054 219922 341122 219978
rect 341178 219922 363250 219978
rect 363306 219922 363374 219978
rect 363430 219922 363498 219978
rect 363554 219922 363622 219978
rect 363678 219922 371718 219978
rect 371774 219922 371842 219978
rect 371898 219922 381250 219978
rect 381306 219922 381374 219978
rect 381430 219922 381498 219978
rect 381554 219922 381622 219978
rect 381678 219922 399250 219978
rect 399306 219922 399374 219978
rect 399430 219922 399498 219978
rect 399554 219922 399622 219978
rect 399678 219922 402438 219978
rect 402494 219922 402562 219978
rect 402618 219922 433158 219978
rect 433214 219922 433282 219978
rect 433338 219922 435250 219978
rect 435306 219922 435374 219978
rect 435430 219922 435498 219978
rect 435554 219922 435622 219978
rect 435678 219922 453250 219978
rect 453306 219922 453374 219978
rect 453430 219922 453498 219978
rect 453554 219922 453622 219978
rect 453678 219922 471250 219978
rect 471306 219922 471374 219978
rect 471430 219922 471498 219978
rect 471554 219922 471622 219978
rect 471678 219922 489250 219978
rect 489306 219922 489374 219978
rect 489430 219922 489498 219978
rect 489554 219922 489622 219978
rect 489678 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 79878 208350
rect 79934 208294 80002 208350
rect 80058 208294 110598 208350
rect 110654 208294 110722 208350
rect 110778 208294 141318 208350
rect 141374 208294 141442 208350
rect 141498 208294 172038 208350
rect 172094 208294 172162 208350
rect 172218 208294 202758 208350
rect 202814 208294 202882 208350
rect 202938 208294 233478 208350
rect 233534 208294 233602 208350
rect 233658 208294 264198 208350
rect 264254 208294 264322 208350
rect 264378 208294 294918 208350
rect 294974 208294 295042 208350
rect 295098 208294 325638 208350
rect 325694 208294 325762 208350
rect 325818 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 356358 208350
rect 356414 208294 356482 208350
rect 356538 208294 366970 208350
rect 367026 208294 367094 208350
rect 367150 208294 367218 208350
rect 367274 208294 367342 208350
rect 367398 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 387078 208350
rect 387134 208294 387202 208350
rect 387258 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 417798 208350
rect 417854 208294 417922 208350
rect 417978 208294 420970 208350
rect 421026 208294 421094 208350
rect 421150 208294 421218 208350
rect 421274 208294 421342 208350
rect 421398 208294 438970 208350
rect 439026 208294 439094 208350
rect 439150 208294 439218 208350
rect 439274 208294 439342 208350
rect 439398 208294 456970 208350
rect 457026 208294 457094 208350
rect 457150 208294 457218 208350
rect 457274 208294 457342 208350
rect 457398 208294 474970 208350
rect 475026 208294 475094 208350
rect 475150 208294 475218 208350
rect 475274 208294 475342 208350
rect 475398 208294 492970 208350
rect 493026 208294 493094 208350
rect 493150 208294 493218 208350
rect 493274 208294 493342 208350
rect 493398 208294 510970 208350
rect 511026 208294 511094 208350
rect 511150 208294 511218 208350
rect 511274 208294 511342 208350
rect 511398 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 79878 208226
rect 79934 208170 80002 208226
rect 80058 208170 110598 208226
rect 110654 208170 110722 208226
rect 110778 208170 141318 208226
rect 141374 208170 141442 208226
rect 141498 208170 172038 208226
rect 172094 208170 172162 208226
rect 172218 208170 202758 208226
rect 202814 208170 202882 208226
rect 202938 208170 233478 208226
rect 233534 208170 233602 208226
rect 233658 208170 264198 208226
rect 264254 208170 264322 208226
rect 264378 208170 294918 208226
rect 294974 208170 295042 208226
rect 295098 208170 325638 208226
rect 325694 208170 325762 208226
rect 325818 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 356358 208226
rect 356414 208170 356482 208226
rect 356538 208170 366970 208226
rect 367026 208170 367094 208226
rect 367150 208170 367218 208226
rect 367274 208170 367342 208226
rect 367398 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 387078 208226
rect 387134 208170 387202 208226
rect 387258 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 417798 208226
rect 417854 208170 417922 208226
rect 417978 208170 420970 208226
rect 421026 208170 421094 208226
rect 421150 208170 421218 208226
rect 421274 208170 421342 208226
rect 421398 208170 438970 208226
rect 439026 208170 439094 208226
rect 439150 208170 439218 208226
rect 439274 208170 439342 208226
rect 439398 208170 456970 208226
rect 457026 208170 457094 208226
rect 457150 208170 457218 208226
rect 457274 208170 457342 208226
rect 457398 208170 474970 208226
rect 475026 208170 475094 208226
rect 475150 208170 475218 208226
rect 475274 208170 475342 208226
rect 475398 208170 492970 208226
rect 493026 208170 493094 208226
rect 493150 208170 493218 208226
rect 493274 208170 493342 208226
rect 493398 208170 510970 208226
rect 511026 208170 511094 208226
rect 511150 208170 511218 208226
rect 511274 208170 511342 208226
rect 511398 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 79878 208102
rect 79934 208046 80002 208102
rect 80058 208046 110598 208102
rect 110654 208046 110722 208102
rect 110778 208046 141318 208102
rect 141374 208046 141442 208102
rect 141498 208046 172038 208102
rect 172094 208046 172162 208102
rect 172218 208046 202758 208102
rect 202814 208046 202882 208102
rect 202938 208046 233478 208102
rect 233534 208046 233602 208102
rect 233658 208046 264198 208102
rect 264254 208046 264322 208102
rect 264378 208046 294918 208102
rect 294974 208046 295042 208102
rect 295098 208046 325638 208102
rect 325694 208046 325762 208102
rect 325818 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 356358 208102
rect 356414 208046 356482 208102
rect 356538 208046 366970 208102
rect 367026 208046 367094 208102
rect 367150 208046 367218 208102
rect 367274 208046 367342 208102
rect 367398 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 387078 208102
rect 387134 208046 387202 208102
rect 387258 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 417798 208102
rect 417854 208046 417922 208102
rect 417978 208046 420970 208102
rect 421026 208046 421094 208102
rect 421150 208046 421218 208102
rect 421274 208046 421342 208102
rect 421398 208046 438970 208102
rect 439026 208046 439094 208102
rect 439150 208046 439218 208102
rect 439274 208046 439342 208102
rect 439398 208046 456970 208102
rect 457026 208046 457094 208102
rect 457150 208046 457218 208102
rect 457274 208046 457342 208102
rect 457398 208046 474970 208102
rect 475026 208046 475094 208102
rect 475150 208046 475218 208102
rect 475274 208046 475342 208102
rect 475398 208046 492970 208102
rect 493026 208046 493094 208102
rect 493150 208046 493218 208102
rect 493274 208046 493342 208102
rect 493398 208046 510970 208102
rect 511026 208046 511094 208102
rect 511150 208046 511218 208102
rect 511274 208046 511342 208102
rect 511398 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 79878 207978
rect 79934 207922 80002 207978
rect 80058 207922 110598 207978
rect 110654 207922 110722 207978
rect 110778 207922 141318 207978
rect 141374 207922 141442 207978
rect 141498 207922 172038 207978
rect 172094 207922 172162 207978
rect 172218 207922 202758 207978
rect 202814 207922 202882 207978
rect 202938 207922 233478 207978
rect 233534 207922 233602 207978
rect 233658 207922 264198 207978
rect 264254 207922 264322 207978
rect 264378 207922 294918 207978
rect 294974 207922 295042 207978
rect 295098 207922 325638 207978
rect 325694 207922 325762 207978
rect 325818 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 356358 207978
rect 356414 207922 356482 207978
rect 356538 207922 366970 207978
rect 367026 207922 367094 207978
rect 367150 207922 367218 207978
rect 367274 207922 367342 207978
rect 367398 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 387078 207978
rect 387134 207922 387202 207978
rect 387258 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 417798 207978
rect 417854 207922 417922 207978
rect 417978 207922 420970 207978
rect 421026 207922 421094 207978
rect 421150 207922 421218 207978
rect 421274 207922 421342 207978
rect 421398 207922 438970 207978
rect 439026 207922 439094 207978
rect 439150 207922 439218 207978
rect 439274 207922 439342 207978
rect 439398 207922 456970 207978
rect 457026 207922 457094 207978
rect 457150 207922 457218 207978
rect 457274 207922 457342 207978
rect 457398 207922 474970 207978
rect 475026 207922 475094 207978
rect 475150 207922 475218 207978
rect 475274 207922 475342 207978
rect 475398 207922 492970 207978
rect 493026 207922 493094 207978
rect 493150 207922 493218 207978
rect 493274 207922 493342 207978
rect 493398 207922 510970 207978
rect 511026 207922 511094 207978
rect 511150 207922 511218 207978
rect 511274 207922 511342 207978
rect 511398 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 64518 202350
rect 64574 202294 64642 202350
rect 64698 202294 95238 202350
rect 95294 202294 95362 202350
rect 95418 202294 125958 202350
rect 126014 202294 126082 202350
rect 126138 202294 156678 202350
rect 156734 202294 156802 202350
rect 156858 202294 187398 202350
rect 187454 202294 187522 202350
rect 187578 202294 218118 202350
rect 218174 202294 218242 202350
rect 218298 202294 248838 202350
rect 248894 202294 248962 202350
rect 249018 202294 279558 202350
rect 279614 202294 279682 202350
rect 279738 202294 310278 202350
rect 310334 202294 310402 202350
rect 310458 202294 340998 202350
rect 341054 202294 341122 202350
rect 341178 202294 363250 202350
rect 363306 202294 363374 202350
rect 363430 202294 363498 202350
rect 363554 202294 363622 202350
rect 363678 202294 371718 202350
rect 371774 202294 371842 202350
rect 371898 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 402438 202350
rect 402494 202294 402562 202350
rect 402618 202294 433158 202350
rect 433214 202294 433282 202350
rect 433338 202294 435250 202350
rect 435306 202294 435374 202350
rect 435430 202294 435498 202350
rect 435554 202294 435622 202350
rect 435678 202294 453250 202350
rect 453306 202294 453374 202350
rect 453430 202294 453498 202350
rect 453554 202294 453622 202350
rect 453678 202294 471250 202350
rect 471306 202294 471374 202350
rect 471430 202294 471498 202350
rect 471554 202294 471622 202350
rect 471678 202294 489250 202350
rect 489306 202294 489374 202350
rect 489430 202294 489498 202350
rect 489554 202294 489622 202350
rect 489678 202294 507250 202350
rect 507306 202294 507374 202350
rect 507430 202294 507498 202350
rect 507554 202294 507622 202350
rect 507678 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 64518 202226
rect 64574 202170 64642 202226
rect 64698 202170 95238 202226
rect 95294 202170 95362 202226
rect 95418 202170 125958 202226
rect 126014 202170 126082 202226
rect 126138 202170 156678 202226
rect 156734 202170 156802 202226
rect 156858 202170 187398 202226
rect 187454 202170 187522 202226
rect 187578 202170 218118 202226
rect 218174 202170 218242 202226
rect 218298 202170 248838 202226
rect 248894 202170 248962 202226
rect 249018 202170 279558 202226
rect 279614 202170 279682 202226
rect 279738 202170 310278 202226
rect 310334 202170 310402 202226
rect 310458 202170 340998 202226
rect 341054 202170 341122 202226
rect 341178 202170 363250 202226
rect 363306 202170 363374 202226
rect 363430 202170 363498 202226
rect 363554 202170 363622 202226
rect 363678 202170 371718 202226
rect 371774 202170 371842 202226
rect 371898 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 402438 202226
rect 402494 202170 402562 202226
rect 402618 202170 433158 202226
rect 433214 202170 433282 202226
rect 433338 202170 435250 202226
rect 435306 202170 435374 202226
rect 435430 202170 435498 202226
rect 435554 202170 435622 202226
rect 435678 202170 453250 202226
rect 453306 202170 453374 202226
rect 453430 202170 453498 202226
rect 453554 202170 453622 202226
rect 453678 202170 471250 202226
rect 471306 202170 471374 202226
rect 471430 202170 471498 202226
rect 471554 202170 471622 202226
rect 471678 202170 489250 202226
rect 489306 202170 489374 202226
rect 489430 202170 489498 202226
rect 489554 202170 489622 202226
rect 489678 202170 507250 202226
rect 507306 202170 507374 202226
rect 507430 202170 507498 202226
rect 507554 202170 507622 202226
rect 507678 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 64518 202102
rect 64574 202046 64642 202102
rect 64698 202046 95238 202102
rect 95294 202046 95362 202102
rect 95418 202046 125958 202102
rect 126014 202046 126082 202102
rect 126138 202046 156678 202102
rect 156734 202046 156802 202102
rect 156858 202046 187398 202102
rect 187454 202046 187522 202102
rect 187578 202046 218118 202102
rect 218174 202046 218242 202102
rect 218298 202046 248838 202102
rect 248894 202046 248962 202102
rect 249018 202046 279558 202102
rect 279614 202046 279682 202102
rect 279738 202046 310278 202102
rect 310334 202046 310402 202102
rect 310458 202046 340998 202102
rect 341054 202046 341122 202102
rect 341178 202046 363250 202102
rect 363306 202046 363374 202102
rect 363430 202046 363498 202102
rect 363554 202046 363622 202102
rect 363678 202046 371718 202102
rect 371774 202046 371842 202102
rect 371898 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 402438 202102
rect 402494 202046 402562 202102
rect 402618 202046 433158 202102
rect 433214 202046 433282 202102
rect 433338 202046 435250 202102
rect 435306 202046 435374 202102
rect 435430 202046 435498 202102
rect 435554 202046 435622 202102
rect 435678 202046 453250 202102
rect 453306 202046 453374 202102
rect 453430 202046 453498 202102
rect 453554 202046 453622 202102
rect 453678 202046 471250 202102
rect 471306 202046 471374 202102
rect 471430 202046 471498 202102
rect 471554 202046 471622 202102
rect 471678 202046 489250 202102
rect 489306 202046 489374 202102
rect 489430 202046 489498 202102
rect 489554 202046 489622 202102
rect 489678 202046 507250 202102
rect 507306 202046 507374 202102
rect 507430 202046 507498 202102
rect 507554 202046 507622 202102
rect 507678 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 64518 201978
rect 64574 201922 64642 201978
rect 64698 201922 95238 201978
rect 95294 201922 95362 201978
rect 95418 201922 125958 201978
rect 126014 201922 126082 201978
rect 126138 201922 156678 201978
rect 156734 201922 156802 201978
rect 156858 201922 187398 201978
rect 187454 201922 187522 201978
rect 187578 201922 218118 201978
rect 218174 201922 218242 201978
rect 218298 201922 248838 201978
rect 248894 201922 248962 201978
rect 249018 201922 279558 201978
rect 279614 201922 279682 201978
rect 279738 201922 310278 201978
rect 310334 201922 310402 201978
rect 310458 201922 340998 201978
rect 341054 201922 341122 201978
rect 341178 201922 363250 201978
rect 363306 201922 363374 201978
rect 363430 201922 363498 201978
rect 363554 201922 363622 201978
rect 363678 201922 371718 201978
rect 371774 201922 371842 201978
rect 371898 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 402438 201978
rect 402494 201922 402562 201978
rect 402618 201922 433158 201978
rect 433214 201922 433282 201978
rect 433338 201922 435250 201978
rect 435306 201922 435374 201978
rect 435430 201922 435498 201978
rect 435554 201922 435622 201978
rect 435678 201922 453250 201978
rect 453306 201922 453374 201978
rect 453430 201922 453498 201978
rect 453554 201922 453622 201978
rect 453678 201922 471250 201978
rect 471306 201922 471374 201978
rect 471430 201922 471498 201978
rect 471554 201922 471622 201978
rect 471678 201922 489250 201978
rect 489306 201922 489374 201978
rect 489430 201922 489498 201978
rect 489554 201922 489622 201978
rect 489678 201922 507250 201978
rect 507306 201922 507374 201978
rect 507430 201922 507498 201978
rect 507554 201922 507622 201978
rect 507678 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 79878 190350
rect 79934 190294 80002 190350
rect 80058 190294 110598 190350
rect 110654 190294 110722 190350
rect 110778 190294 141318 190350
rect 141374 190294 141442 190350
rect 141498 190294 172038 190350
rect 172094 190294 172162 190350
rect 172218 190294 202758 190350
rect 202814 190294 202882 190350
rect 202938 190294 233478 190350
rect 233534 190294 233602 190350
rect 233658 190294 264198 190350
rect 264254 190294 264322 190350
rect 264378 190294 294918 190350
rect 294974 190294 295042 190350
rect 295098 190294 325638 190350
rect 325694 190294 325762 190350
rect 325818 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 356358 190350
rect 356414 190294 356482 190350
rect 356538 190294 366970 190350
rect 367026 190294 367094 190350
rect 367150 190294 367218 190350
rect 367274 190294 367342 190350
rect 367398 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 387078 190350
rect 387134 190294 387202 190350
rect 387258 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 417798 190350
rect 417854 190294 417922 190350
rect 417978 190294 420970 190350
rect 421026 190294 421094 190350
rect 421150 190294 421218 190350
rect 421274 190294 421342 190350
rect 421398 190294 438970 190350
rect 439026 190294 439094 190350
rect 439150 190294 439218 190350
rect 439274 190294 439342 190350
rect 439398 190294 456970 190350
rect 457026 190294 457094 190350
rect 457150 190294 457218 190350
rect 457274 190294 457342 190350
rect 457398 190294 474970 190350
rect 475026 190294 475094 190350
rect 475150 190294 475218 190350
rect 475274 190294 475342 190350
rect 475398 190294 492970 190350
rect 493026 190294 493094 190350
rect 493150 190294 493218 190350
rect 493274 190294 493342 190350
rect 493398 190294 510970 190350
rect 511026 190294 511094 190350
rect 511150 190294 511218 190350
rect 511274 190294 511342 190350
rect 511398 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 79878 190226
rect 79934 190170 80002 190226
rect 80058 190170 110598 190226
rect 110654 190170 110722 190226
rect 110778 190170 141318 190226
rect 141374 190170 141442 190226
rect 141498 190170 172038 190226
rect 172094 190170 172162 190226
rect 172218 190170 202758 190226
rect 202814 190170 202882 190226
rect 202938 190170 233478 190226
rect 233534 190170 233602 190226
rect 233658 190170 264198 190226
rect 264254 190170 264322 190226
rect 264378 190170 294918 190226
rect 294974 190170 295042 190226
rect 295098 190170 325638 190226
rect 325694 190170 325762 190226
rect 325818 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 356358 190226
rect 356414 190170 356482 190226
rect 356538 190170 366970 190226
rect 367026 190170 367094 190226
rect 367150 190170 367218 190226
rect 367274 190170 367342 190226
rect 367398 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 387078 190226
rect 387134 190170 387202 190226
rect 387258 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 417798 190226
rect 417854 190170 417922 190226
rect 417978 190170 420970 190226
rect 421026 190170 421094 190226
rect 421150 190170 421218 190226
rect 421274 190170 421342 190226
rect 421398 190170 438970 190226
rect 439026 190170 439094 190226
rect 439150 190170 439218 190226
rect 439274 190170 439342 190226
rect 439398 190170 456970 190226
rect 457026 190170 457094 190226
rect 457150 190170 457218 190226
rect 457274 190170 457342 190226
rect 457398 190170 474970 190226
rect 475026 190170 475094 190226
rect 475150 190170 475218 190226
rect 475274 190170 475342 190226
rect 475398 190170 492970 190226
rect 493026 190170 493094 190226
rect 493150 190170 493218 190226
rect 493274 190170 493342 190226
rect 493398 190170 510970 190226
rect 511026 190170 511094 190226
rect 511150 190170 511218 190226
rect 511274 190170 511342 190226
rect 511398 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 79878 190102
rect 79934 190046 80002 190102
rect 80058 190046 110598 190102
rect 110654 190046 110722 190102
rect 110778 190046 141318 190102
rect 141374 190046 141442 190102
rect 141498 190046 172038 190102
rect 172094 190046 172162 190102
rect 172218 190046 202758 190102
rect 202814 190046 202882 190102
rect 202938 190046 233478 190102
rect 233534 190046 233602 190102
rect 233658 190046 264198 190102
rect 264254 190046 264322 190102
rect 264378 190046 294918 190102
rect 294974 190046 295042 190102
rect 295098 190046 325638 190102
rect 325694 190046 325762 190102
rect 325818 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 356358 190102
rect 356414 190046 356482 190102
rect 356538 190046 366970 190102
rect 367026 190046 367094 190102
rect 367150 190046 367218 190102
rect 367274 190046 367342 190102
rect 367398 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 387078 190102
rect 387134 190046 387202 190102
rect 387258 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 417798 190102
rect 417854 190046 417922 190102
rect 417978 190046 420970 190102
rect 421026 190046 421094 190102
rect 421150 190046 421218 190102
rect 421274 190046 421342 190102
rect 421398 190046 438970 190102
rect 439026 190046 439094 190102
rect 439150 190046 439218 190102
rect 439274 190046 439342 190102
rect 439398 190046 456970 190102
rect 457026 190046 457094 190102
rect 457150 190046 457218 190102
rect 457274 190046 457342 190102
rect 457398 190046 474970 190102
rect 475026 190046 475094 190102
rect 475150 190046 475218 190102
rect 475274 190046 475342 190102
rect 475398 190046 492970 190102
rect 493026 190046 493094 190102
rect 493150 190046 493218 190102
rect 493274 190046 493342 190102
rect 493398 190046 510970 190102
rect 511026 190046 511094 190102
rect 511150 190046 511218 190102
rect 511274 190046 511342 190102
rect 511398 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 79878 189978
rect 79934 189922 80002 189978
rect 80058 189922 110598 189978
rect 110654 189922 110722 189978
rect 110778 189922 141318 189978
rect 141374 189922 141442 189978
rect 141498 189922 172038 189978
rect 172094 189922 172162 189978
rect 172218 189922 202758 189978
rect 202814 189922 202882 189978
rect 202938 189922 233478 189978
rect 233534 189922 233602 189978
rect 233658 189922 264198 189978
rect 264254 189922 264322 189978
rect 264378 189922 294918 189978
rect 294974 189922 295042 189978
rect 295098 189922 325638 189978
rect 325694 189922 325762 189978
rect 325818 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 356358 189978
rect 356414 189922 356482 189978
rect 356538 189922 366970 189978
rect 367026 189922 367094 189978
rect 367150 189922 367218 189978
rect 367274 189922 367342 189978
rect 367398 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 387078 189978
rect 387134 189922 387202 189978
rect 387258 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 417798 189978
rect 417854 189922 417922 189978
rect 417978 189922 420970 189978
rect 421026 189922 421094 189978
rect 421150 189922 421218 189978
rect 421274 189922 421342 189978
rect 421398 189922 438970 189978
rect 439026 189922 439094 189978
rect 439150 189922 439218 189978
rect 439274 189922 439342 189978
rect 439398 189922 456970 189978
rect 457026 189922 457094 189978
rect 457150 189922 457218 189978
rect 457274 189922 457342 189978
rect 457398 189922 474970 189978
rect 475026 189922 475094 189978
rect 475150 189922 475218 189978
rect 475274 189922 475342 189978
rect 475398 189922 492970 189978
rect 493026 189922 493094 189978
rect 493150 189922 493218 189978
rect 493274 189922 493342 189978
rect 493398 189922 510970 189978
rect 511026 189922 511094 189978
rect 511150 189922 511218 189978
rect 511274 189922 511342 189978
rect 511398 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 64518 184350
rect 64574 184294 64642 184350
rect 64698 184294 95238 184350
rect 95294 184294 95362 184350
rect 95418 184294 125958 184350
rect 126014 184294 126082 184350
rect 126138 184294 156678 184350
rect 156734 184294 156802 184350
rect 156858 184294 187398 184350
rect 187454 184294 187522 184350
rect 187578 184294 218118 184350
rect 218174 184294 218242 184350
rect 218298 184294 248838 184350
rect 248894 184294 248962 184350
rect 249018 184294 279558 184350
rect 279614 184294 279682 184350
rect 279738 184294 310278 184350
rect 310334 184294 310402 184350
rect 310458 184294 340998 184350
rect 341054 184294 341122 184350
rect 341178 184294 363250 184350
rect 363306 184294 363374 184350
rect 363430 184294 363498 184350
rect 363554 184294 363622 184350
rect 363678 184294 371718 184350
rect 371774 184294 371842 184350
rect 371898 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 402438 184350
rect 402494 184294 402562 184350
rect 402618 184294 433158 184350
rect 433214 184294 433282 184350
rect 433338 184294 435250 184350
rect 435306 184294 435374 184350
rect 435430 184294 435498 184350
rect 435554 184294 435622 184350
rect 435678 184294 453250 184350
rect 453306 184294 453374 184350
rect 453430 184294 453498 184350
rect 453554 184294 453622 184350
rect 453678 184294 471250 184350
rect 471306 184294 471374 184350
rect 471430 184294 471498 184350
rect 471554 184294 471622 184350
rect 471678 184294 489250 184350
rect 489306 184294 489374 184350
rect 489430 184294 489498 184350
rect 489554 184294 489622 184350
rect 489678 184294 507250 184350
rect 507306 184294 507374 184350
rect 507430 184294 507498 184350
rect 507554 184294 507622 184350
rect 507678 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 64518 184226
rect 64574 184170 64642 184226
rect 64698 184170 95238 184226
rect 95294 184170 95362 184226
rect 95418 184170 125958 184226
rect 126014 184170 126082 184226
rect 126138 184170 156678 184226
rect 156734 184170 156802 184226
rect 156858 184170 187398 184226
rect 187454 184170 187522 184226
rect 187578 184170 218118 184226
rect 218174 184170 218242 184226
rect 218298 184170 248838 184226
rect 248894 184170 248962 184226
rect 249018 184170 279558 184226
rect 279614 184170 279682 184226
rect 279738 184170 310278 184226
rect 310334 184170 310402 184226
rect 310458 184170 340998 184226
rect 341054 184170 341122 184226
rect 341178 184170 363250 184226
rect 363306 184170 363374 184226
rect 363430 184170 363498 184226
rect 363554 184170 363622 184226
rect 363678 184170 371718 184226
rect 371774 184170 371842 184226
rect 371898 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 402438 184226
rect 402494 184170 402562 184226
rect 402618 184170 433158 184226
rect 433214 184170 433282 184226
rect 433338 184170 435250 184226
rect 435306 184170 435374 184226
rect 435430 184170 435498 184226
rect 435554 184170 435622 184226
rect 435678 184170 453250 184226
rect 453306 184170 453374 184226
rect 453430 184170 453498 184226
rect 453554 184170 453622 184226
rect 453678 184170 471250 184226
rect 471306 184170 471374 184226
rect 471430 184170 471498 184226
rect 471554 184170 471622 184226
rect 471678 184170 489250 184226
rect 489306 184170 489374 184226
rect 489430 184170 489498 184226
rect 489554 184170 489622 184226
rect 489678 184170 507250 184226
rect 507306 184170 507374 184226
rect 507430 184170 507498 184226
rect 507554 184170 507622 184226
rect 507678 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 64518 184102
rect 64574 184046 64642 184102
rect 64698 184046 95238 184102
rect 95294 184046 95362 184102
rect 95418 184046 125958 184102
rect 126014 184046 126082 184102
rect 126138 184046 156678 184102
rect 156734 184046 156802 184102
rect 156858 184046 187398 184102
rect 187454 184046 187522 184102
rect 187578 184046 218118 184102
rect 218174 184046 218242 184102
rect 218298 184046 248838 184102
rect 248894 184046 248962 184102
rect 249018 184046 279558 184102
rect 279614 184046 279682 184102
rect 279738 184046 310278 184102
rect 310334 184046 310402 184102
rect 310458 184046 340998 184102
rect 341054 184046 341122 184102
rect 341178 184046 363250 184102
rect 363306 184046 363374 184102
rect 363430 184046 363498 184102
rect 363554 184046 363622 184102
rect 363678 184046 371718 184102
rect 371774 184046 371842 184102
rect 371898 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 402438 184102
rect 402494 184046 402562 184102
rect 402618 184046 433158 184102
rect 433214 184046 433282 184102
rect 433338 184046 435250 184102
rect 435306 184046 435374 184102
rect 435430 184046 435498 184102
rect 435554 184046 435622 184102
rect 435678 184046 453250 184102
rect 453306 184046 453374 184102
rect 453430 184046 453498 184102
rect 453554 184046 453622 184102
rect 453678 184046 471250 184102
rect 471306 184046 471374 184102
rect 471430 184046 471498 184102
rect 471554 184046 471622 184102
rect 471678 184046 489250 184102
rect 489306 184046 489374 184102
rect 489430 184046 489498 184102
rect 489554 184046 489622 184102
rect 489678 184046 507250 184102
rect 507306 184046 507374 184102
rect 507430 184046 507498 184102
rect 507554 184046 507622 184102
rect 507678 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 64518 183978
rect 64574 183922 64642 183978
rect 64698 183922 95238 183978
rect 95294 183922 95362 183978
rect 95418 183922 125958 183978
rect 126014 183922 126082 183978
rect 126138 183922 156678 183978
rect 156734 183922 156802 183978
rect 156858 183922 187398 183978
rect 187454 183922 187522 183978
rect 187578 183922 218118 183978
rect 218174 183922 218242 183978
rect 218298 183922 248838 183978
rect 248894 183922 248962 183978
rect 249018 183922 279558 183978
rect 279614 183922 279682 183978
rect 279738 183922 310278 183978
rect 310334 183922 310402 183978
rect 310458 183922 340998 183978
rect 341054 183922 341122 183978
rect 341178 183922 363250 183978
rect 363306 183922 363374 183978
rect 363430 183922 363498 183978
rect 363554 183922 363622 183978
rect 363678 183922 371718 183978
rect 371774 183922 371842 183978
rect 371898 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 402438 183978
rect 402494 183922 402562 183978
rect 402618 183922 433158 183978
rect 433214 183922 433282 183978
rect 433338 183922 435250 183978
rect 435306 183922 435374 183978
rect 435430 183922 435498 183978
rect 435554 183922 435622 183978
rect 435678 183922 453250 183978
rect 453306 183922 453374 183978
rect 453430 183922 453498 183978
rect 453554 183922 453622 183978
rect 453678 183922 471250 183978
rect 471306 183922 471374 183978
rect 471430 183922 471498 183978
rect 471554 183922 471622 183978
rect 471678 183922 489250 183978
rect 489306 183922 489374 183978
rect 489430 183922 489498 183978
rect 489554 183922 489622 183978
rect 489678 183922 507250 183978
rect 507306 183922 507374 183978
rect 507430 183922 507498 183978
rect 507554 183922 507622 183978
rect 507678 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 79878 172350
rect 79934 172294 80002 172350
rect 80058 172294 110598 172350
rect 110654 172294 110722 172350
rect 110778 172294 141318 172350
rect 141374 172294 141442 172350
rect 141498 172294 172038 172350
rect 172094 172294 172162 172350
rect 172218 172294 202758 172350
rect 202814 172294 202882 172350
rect 202938 172294 233478 172350
rect 233534 172294 233602 172350
rect 233658 172294 264198 172350
rect 264254 172294 264322 172350
rect 264378 172294 294918 172350
rect 294974 172294 295042 172350
rect 295098 172294 325638 172350
rect 325694 172294 325762 172350
rect 325818 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 356358 172350
rect 356414 172294 356482 172350
rect 356538 172294 366970 172350
rect 367026 172294 367094 172350
rect 367150 172294 367218 172350
rect 367274 172294 367342 172350
rect 367398 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 387078 172350
rect 387134 172294 387202 172350
rect 387258 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 417798 172350
rect 417854 172294 417922 172350
rect 417978 172294 420970 172350
rect 421026 172294 421094 172350
rect 421150 172294 421218 172350
rect 421274 172294 421342 172350
rect 421398 172294 438970 172350
rect 439026 172294 439094 172350
rect 439150 172294 439218 172350
rect 439274 172294 439342 172350
rect 439398 172294 456970 172350
rect 457026 172294 457094 172350
rect 457150 172294 457218 172350
rect 457274 172294 457342 172350
rect 457398 172294 474970 172350
rect 475026 172294 475094 172350
rect 475150 172294 475218 172350
rect 475274 172294 475342 172350
rect 475398 172294 492970 172350
rect 493026 172294 493094 172350
rect 493150 172294 493218 172350
rect 493274 172294 493342 172350
rect 493398 172294 510970 172350
rect 511026 172294 511094 172350
rect 511150 172294 511218 172350
rect 511274 172294 511342 172350
rect 511398 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 79878 172226
rect 79934 172170 80002 172226
rect 80058 172170 110598 172226
rect 110654 172170 110722 172226
rect 110778 172170 141318 172226
rect 141374 172170 141442 172226
rect 141498 172170 172038 172226
rect 172094 172170 172162 172226
rect 172218 172170 202758 172226
rect 202814 172170 202882 172226
rect 202938 172170 233478 172226
rect 233534 172170 233602 172226
rect 233658 172170 264198 172226
rect 264254 172170 264322 172226
rect 264378 172170 294918 172226
rect 294974 172170 295042 172226
rect 295098 172170 325638 172226
rect 325694 172170 325762 172226
rect 325818 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 356358 172226
rect 356414 172170 356482 172226
rect 356538 172170 366970 172226
rect 367026 172170 367094 172226
rect 367150 172170 367218 172226
rect 367274 172170 367342 172226
rect 367398 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 387078 172226
rect 387134 172170 387202 172226
rect 387258 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 417798 172226
rect 417854 172170 417922 172226
rect 417978 172170 420970 172226
rect 421026 172170 421094 172226
rect 421150 172170 421218 172226
rect 421274 172170 421342 172226
rect 421398 172170 438970 172226
rect 439026 172170 439094 172226
rect 439150 172170 439218 172226
rect 439274 172170 439342 172226
rect 439398 172170 456970 172226
rect 457026 172170 457094 172226
rect 457150 172170 457218 172226
rect 457274 172170 457342 172226
rect 457398 172170 474970 172226
rect 475026 172170 475094 172226
rect 475150 172170 475218 172226
rect 475274 172170 475342 172226
rect 475398 172170 492970 172226
rect 493026 172170 493094 172226
rect 493150 172170 493218 172226
rect 493274 172170 493342 172226
rect 493398 172170 510970 172226
rect 511026 172170 511094 172226
rect 511150 172170 511218 172226
rect 511274 172170 511342 172226
rect 511398 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 79878 172102
rect 79934 172046 80002 172102
rect 80058 172046 110598 172102
rect 110654 172046 110722 172102
rect 110778 172046 141318 172102
rect 141374 172046 141442 172102
rect 141498 172046 172038 172102
rect 172094 172046 172162 172102
rect 172218 172046 202758 172102
rect 202814 172046 202882 172102
rect 202938 172046 233478 172102
rect 233534 172046 233602 172102
rect 233658 172046 264198 172102
rect 264254 172046 264322 172102
rect 264378 172046 294918 172102
rect 294974 172046 295042 172102
rect 295098 172046 325638 172102
rect 325694 172046 325762 172102
rect 325818 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 356358 172102
rect 356414 172046 356482 172102
rect 356538 172046 366970 172102
rect 367026 172046 367094 172102
rect 367150 172046 367218 172102
rect 367274 172046 367342 172102
rect 367398 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 387078 172102
rect 387134 172046 387202 172102
rect 387258 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 417798 172102
rect 417854 172046 417922 172102
rect 417978 172046 420970 172102
rect 421026 172046 421094 172102
rect 421150 172046 421218 172102
rect 421274 172046 421342 172102
rect 421398 172046 438970 172102
rect 439026 172046 439094 172102
rect 439150 172046 439218 172102
rect 439274 172046 439342 172102
rect 439398 172046 456970 172102
rect 457026 172046 457094 172102
rect 457150 172046 457218 172102
rect 457274 172046 457342 172102
rect 457398 172046 474970 172102
rect 475026 172046 475094 172102
rect 475150 172046 475218 172102
rect 475274 172046 475342 172102
rect 475398 172046 492970 172102
rect 493026 172046 493094 172102
rect 493150 172046 493218 172102
rect 493274 172046 493342 172102
rect 493398 172046 510970 172102
rect 511026 172046 511094 172102
rect 511150 172046 511218 172102
rect 511274 172046 511342 172102
rect 511398 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 79878 171978
rect 79934 171922 80002 171978
rect 80058 171922 110598 171978
rect 110654 171922 110722 171978
rect 110778 171922 141318 171978
rect 141374 171922 141442 171978
rect 141498 171922 172038 171978
rect 172094 171922 172162 171978
rect 172218 171922 202758 171978
rect 202814 171922 202882 171978
rect 202938 171922 233478 171978
rect 233534 171922 233602 171978
rect 233658 171922 264198 171978
rect 264254 171922 264322 171978
rect 264378 171922 294918 171978
rect 294974 171922 295042 171978
rect 295098 171922 325638 171978
rect 325694 171922 325762 171978
rect 325818 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 356358 171978
rect 356414 171922 356482 171978
rect 356538 171922 366970 171978
rect 367026 171922 367094 171978
rect 367150 171922 367218 171978
rect 367274 171922 367342 171978
rect 367398 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 387078 171978
rect 387134 171922 387202 171978
rect 387258 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 417798 171978
rect 417854 171922 417922 171978
rect 417978 171922 420970 171978
rect 421026 171922 421094 171978
rect 421150 171922 421218 171978
rect 421274 171922 421342 171978
rect 421398 171922 438970 171978
rect 439026 171922 439094 171978
rect 439150 171922 439218 171978
rect 439274 171922 439342 171978
rect 439398 171922 456970 171978
rect 457026 171922 457094 171978
rect 457150 171922 457218 171978
rect 457274 171922 457342 171978
rect 457398 171922 474970 171978
rect 475026 171922 475094 171978
rect 475150 171922 475218 171978
rect 475274 171922 475342 171978
rect 475398 171922 492970 171978
rect 493026 171922 493094 171978
rect 493150 171922 493218 171978
rect 493274 171922 493342 171978
rect 493398 171922 510970 171978
rect 511026 171922 511094 171978
rect 511150 171922 511218 171978
rect 511274 171922 511342 171978
rect 511398 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 64518 166350
rect 64574 166294 64642 166350
rect 64698 166294 95238 166350
rect 95294 166294 95362 166350
rect 95418 166294 125958 166350
rect 126014 166294 126082 166350
rect 126138 166294 156678 166350
rect 156734 166294 156802 166350
rect 156858 166294 187398 166350
rect 187454 166294 187522 166350
rect 187578 166294 218118 166350
rect 218174 166294 218242 166350
rect 218298 166294 248838 166350
rect 248894 166294 248962 166350
rect 249018 166294 279558 166350
rect 279614 166294 279682 166350
rect 279738 166294 310278 166350
rect 310334 166294 310402 166350
rect 310458 166294 340998 166350
rect 341054 166294 341122 166350
rect 341178 166294 363250 166350
rect 363306 166294 363374 166350
rect 363430 166294 363498 166350
rect 363554 166294 363622 166350
rect 363678 166294 371718 166350
rect 371774 166294 371842 166350
rect 371898 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 402438 166350
rect 402494 166294 402562 166350
rect 402618 166294 433158 166350
rect 433214 166294 433282 166350
rect 433338 166294 435250 166350
rect 435306 166294 435374 166350
rect 435430 166294 435498 166350
rect 435554 166294 435622 166350
rect 435678 166294 453250 166350
rect 453306 166294 453374 166350
rect 453430 166294 453498 166350
rect 453554 166294 453622 166350
rect 453678 166294 471250 166350
rect 471306 166294 471374 166350
rect 471430 166294 471498 166350
rect 471554 166294 471622 166350
rect 471678 166294 489250 166350
rect 489306 166294 489374 166350
rect 489430 166294 489498 166350
rect 489554 166294 489622 166350
rect 489678 166294 507250 166350
rect 507306 166294 507374 166350
rect 507430 166294 507498 166350
rect 507554 166294 507622 166350
rect 507678 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 64518 166226
rect 64574 166170 64642 166226
rect 64698 166170 95238 166226
rect 95294 166170 95362 166226
rect 95418 166170 125958 166226
rect 126014 166170 126082 166226
rect 126138 166170 156678 166226
rect 156734 166170 156802 166226
rect 156858 166170 187398 166226
rect 187454 166170 187522 166226
rect 187578 166170 218118 166226
rect 218174 166170 218242 166226
rect 218298 166170 248838 166226
rect 248894 166170 248962 166226
rect 249018 166170 279558 166226
rect 279614 166170 279682 166226
rect 279738 166170 310278 166226
rect 310334 166170 310402 166226
rect 310458 166170 340998 166226
rect 341054 166170 341122 166226
rect 341178 166170 363250 166226
rect 363306 166170 363374 166226
rect 363430 166170 363498 166226
rect 363554 166170 363622 166226
rect 363678 166170 371718 166226
rect 371774 166170 371842 166226
rect 371898 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 402438 166226
rect 402494 166170 402562 166226
rect 402618 166170 433158 166226
rect 433214 166170 433282 166226
rect 433338 166170 435250 166226
rect 435306 166170 435374 166226
rect 435430 166170 435498 166226
rect 435554 166170 435622 166226
rect 435678 166170 453250 166226
rect 453306 166170 453374 166226
rect 453430 166170 453498 166226
rect 453554 166170 453622 166226
rect 453678 166170 471250 166226
rect 471306 166170 471374 166226
rect 471430 166170 471498 166226
rect 471554 166170 471622 166226
rect 471678 166170 489250 166226
rect 489306 166170 489374 166226
rect 489430 166170 489498 166226
rect 489554 166170 489622 166226
rect 489678 166170 507250 166226
rect 507306 166170 507374 166226
rect 507430 166170 507498 166226
rect 507554 166170 507622 166226
rect 507678 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 64518 166102
rect 64574 166046 64642 166102
rect 64698 166046 95238 166102
rect 95294 166046 95362 166102
rect 95418 166046 125958 166102
rect 126014 166046 126082 166102
rect 126138 166046 156678 166102
rect 156734 166046 156802 166102
rect 156858 166046 187398 166102
rect 187454 166046 187522 166102
rect 187578 166046 218118 166102
rect 218174 166046 218242 166102
rect 218298 166046 248838 166102
rect 248894 166046 248962 166102
rect 249018 166046 279558 166102
rect 279614 166046 279682 166102
rect 279738 166046 310278 166102
rect 310334 166046 310402 166102
rect 310458 166046 340998 166102
rect 341054 166046 341122 166102
rect 341178 166046 363250 166102
rect 363306 166046 363374 166102
rect 363430 166046 363498 166102
rect 363554 166046 363622 166102
rect 363678 166046 371718 166102
rect 371774 166046 371842 166102
rect 371898 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 402438 166102
rect 402494 166046 402562 166102
rect 402618 166046 433158 166102
rect 433214 166046 433282 166102
rect 433338 166046 435250 166102
rect 435306 166046 435374 166102
rect 435430 166046 435498 166102
rect 435554 166046 435622 166102
rect 435678 166046 453250 166102
rect 453306 166046 453374 166102
rect 453430 166046 453498 166102
rect 453554 166046 453622 166102
rect 453678 166046 471250 166102
rect 471306 166046 471374 166102
rect 471430 166046 471498 166102
rect 471554 166046 471622 166102
rect 471678 166046 489250 166102
rect 489306 166046 489374 166102
rect 489430 166046 489498 166102
rect 489554 166046 489622 166102
rect 489678 166046 507250 166102
rect 507306 166046 507374 166102
rect 507430 166046 507498 166102
rect 507554 166046 507622 166102
rect 507678 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 64518 165978
rect 64574 165922 64642 165978
rect 64698 165922 95238 165978
rect 95294 165922 95362 165978
rect 95418 165922 125958 165978
rect 126014 165922 126082 165978
rect 126138 165922 156678 165978
rect 156734 165922 156802 165978
rect 156858 165922 187398 165978
rect 187454 165922 187522 165978
rect 187578 165922 218118 165978
rect 218174 165922 218242 165978
rect 218298 165922 248838 165978
rect 248894 165922 248962 165978
rect 249018 165922 279558 165978
rect 279614 165922 279682 165978
rect 279738 165922 310278 165978
rect 310334 165922 310402 165978
rect 310458 165922 340998 165978
rect 341054 165922 341122 165978
rect 341178 165922 363250 165978
rect 363306 165922 363374 165978
rect 363430 165922 363498 165978
rect 363554 165922 363622 165978
rect 363678 165922 371718 165978
rect 371774 165922 371842 165978
rect 371898 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 402438 165978
rect 402494 165922 402562 165978
rect 402618 165922 433158 165978
rect 433214 165922 433282 165978
rect 433338 165922 435250 165978
rect 435306 165922 435374 165978
rect 435430 165922 435498 165978
rect 435554 165922 435622 165978
rect 435678 165922 453250 165978
rect 453306 165922 453374 165978
rect 453430 165922 453498 165978
rect 453554 165922 453622 165978
rect 453678 165922 471250 165978
rect 471306 165922 471374 165978
rect 471430 165922 471498 165978
rect 471554 165922 471622 165978
rect 471678 165922 489250 165978
rect 489306 165922 489374 165978
rect 489430 165922 489498 165978
rect 489554 165922 489622 165978
rect 489678 165922 507250 165978
rect 507306 165922 507374 165978
rect 507430 165922 507498 165978
rect 507554 165922 507622 165978
rect 507678 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 79878 154350
rect 79934 154294 80002 154350
rect 80058 154294 110598 154350
rect 110654 154294 110722 154350
rect 110778 154294 141318 154350
rect 141374 154294 141442 154350
rect 141498 154294 172038 154350
rect 172094 154294 172162 154350
rect 172218 154294 202758 154350
rect 202814 154294 202882 154350
rect 202938 154294 233478 154350
rect 233534 154294 233602 154350
rect 233658 154294 264198 154350
rect 264254 154294 264322 154350
rect 264378 154294 294918 154350
rect 294974 154294 295042 154350
rect 295098 154294 325638 154350
rect 325694 154294 325762 154350
rect 325818 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 356358 154350
rect 356414 154294 356482 154350
rect 356538 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 387078 154350
rect 387134 154294 387202 154350
rect 387258 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 417798 154350
rect 417854 154294 417922 154350
rect 417978 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 79878 154226
rect 79934 154170 80002 154226
rect 80058 154170 110598 154226
rect 110654 154170 110722 154226
rect 110778 154170 141318 154226
rect 141374 154170 141442 154226
rect 141498 154170 172038 154226
rect 172094 154170 172162 154226
rect 172218 154170 202758 154226
rect 202814 154170 202882 154226
rect 202938 154170 233478 154226
rect 233534 154170 233602 154226
rect 233658 154170 264198 154226
rect 264254 154170 264322 154226
rect 264378 154170 294918 154226
rect 294974 154170 295042 154226
rect 295098 154170 325638 154226
rect 325694 154170 325762 154226
rect 325818 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 356358 154226
rect 356414 154170 356482 154226
rect 356538 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 387078 154226
rect 387134 154170 387202 154226
rect 387258 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 417798 154226
rect 417854 154170 417922 154226
rect 417978 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 79878 154102
rect 79934 154046 80002 154102
rect 80058 154046 110598 154102
rect 110654 154046 110722 154102
rect 110778 154046 141318 154102
rect 141374 154046 141442 154102
rect 141498 154046 172038 154102
rect 172094 154046 172162 154102
rect 172218 154046 202758 154102
rect 202814 154046 202882 154102
rect 202938 154046 233478 154102
rect 233534 154046 233602 154102
rect 233658 154046 264198 154102
rect 264254 154046 264322 154102
rect 264378 154046 294918 154102
rect 294974 154046 295042 154102
rect 295098 154046 325638 154102
rect 325694 154046 325762 154102
rect 325818 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 356358 154102
rect 356414 154046 356482 154102
rect 356538 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 387078 154102
rect 387134 154046 387202 154102
rect 387258 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 417798 154102
rect 417854 154046 417922 154102
rect 417978 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 79878 153978
rect 79934 153922 80002 153978
rect 80058 153922 110598 153978
rect 110654 153922 110722 153978
rect 110778 153922 141318 153978
rect 141374 153922 141442 153978
rect 141498 153922 172038 153978
rect 172094 153922 172162 153978
rect 172218 153922 202758 153978
rect 202814 153922 202882 153978
rect 202938 153922 233478 153978
rect 233534 153922 233602 153978
rect 233658 153922 264198 153978
rect 264254 153922 264322 153978
rect 264378 153922 294918 153978
rect 294974 153922 295042 153978
rect 295098 153922 325638 153978
rect 325694 153922 325762 153978
rect 325818 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 356358 153978
rect 356414 153922 356482 153978
rect 356538 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 387078 153978
rect 387134 153922 387202 153978
rect 387258 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 417798 153978
rect 417854 153922 417922 153978
rect 417978 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 64518 148350
rect 64574 148294 64642 148350
rect 64698 148294 95238 148350
rect 95294 148294 95362 148350
rect 95418 148294 125958 148350
rect 126014 148294 126082 148350
rect 126138 148294 156678 148350
rect 156734 148294 156802 148350
rect 156858 148294 187398 148350
rect 187454 148294 187522 148350
rect 187578 148294 218118 148350
rect 218174 148294 218242 148350
rect 218298 148294 248838 148350
rect 248894 148294 248962 148350
rect 249018 148294 279558 148350
rect 279614 148294 279682 148350
rect 279738 148294 310278 148350
rect 310334 148294 310402 148350
rect 310458 148294 340998 148350
rect 341054 148294 341122 148350
rect 341178 148294 363250 148350
rect 363306 148294 363374 148350
rect 363430 148294 363498 148350
rect 363554 148294 363622 148350
rect 363678 148294 371718 148350
rect 371774 148294 371842 148350
rect 371898 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 402438 148350
rect 402494 148294 402562 148350
rect 402618 148294 433158 148350
rect 433214 148294 433282 148350
rect 433338 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 64518 148226
rect 64574 148170 64642 148226
rect 64698 148170 95238 148226
rect 95294 148170 95362 148226
rect 95418 148170 125958 148226
rect 126014 148170 126082 148226
rect 126138 148170 156678 148226
rect 156734 148170 156802 148226
rect 156858 148170 187398 148226
rect 187454 148170 187522 148226
rect 187578 148170 218118 148226
rect 218174 148170 218242 148226
rect 218298 148170 248838 148226
rect 248894 148170 248962 148226
rect 249018 148170 279558 148226
rect 279614 148170 279682 148226
rect 279738 148170 310278 148226
rect 310334 148170 310402 148226
rect 310458 148170 340998 148226
rect 341054 148170 341122 148226
rect 341178 148170 363250 148226
rect 363306 148170 363374 148226
rect 363430 148170 363498 148226
rect 363554 148170 363622 148226
rect 363678 148170 371718 148226
rect 371774 148170 371842 148226
rect 371898 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 402438 148226
rect 402494 148170 402562 148226
rect 402618 148170 433158 148226
rect 433214 148170 433282 148226
rect 433338 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 64518 148102
rect 64574 148046 64642 148102
rect 64698 148046 95238 148102
rect 95294 148046 95362 148102
rect 95418 148046 125958 148102
rect 126014 148046 126082 148102
rect 126138 148046 156678 148102
rect 156734 148046 156802 148102
rect 156858 148046 187398 148102
rect 187454 148046 187522 148102
rect 187578 148046 218118 148102
rect 218174 148046 218242 148102
rect 218298 148046 248838 148102
rect 248894 148046 248962 148102
rect 249018 148046 279558 148102
rect 279614 148046 279682 148102
rect 279738 148046 310278 148102
rect 310334 148046 310402 148102
rect 310458 148046 340998 148102
rect 341054 148046 341122 148102
rect 341178 148046 363250 148102
rect 363306 148046 363374 148102
rect 363430 148046 363498 148102
rect 363554 148046 363622 148102
rect 363678 148046 371718 148102
rect 371774 148046 371842 148102
rect 371898 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 402438 148102
rect 402494 148046 402562 148102
rect 402618 148046 433158 148102
rect 433214 148046 433282 148102
rect 433338 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 64518 147978
rect 64574 147922 64642 147978
rect 64698 147922 95238 147978
rect 95294 147922 95362 147978
rect 95418 147922 125958 147978
rect 126014 147922 126082 147978
rect 126138 147922 156678 147978
rect 156734 147922 156802 147978
rect 156858 147922 187398 147978
rect 187454 147922 187522 147978
rect 187578 147922 218118 147978
rect 218174 147922 218242 147978
rect 218298 147922 248838 147978
rect 248894 147922 248962 147978
rect 249018 147922 279558 147978
rect 279614 147922 279682 147978
rect 279738 147922 310278 147978
rect 310334 147922 310402 147978
rect 310458 147922 340998 147978
rect 341054 147922 341122 147978
rect 341178 147922 363250 147978
rect 363306 147922 363374 147978
rect 363430 147922 363498 147978
rect 363554 147922 363622 147978
rect 363678 147922 371718 147978
rect 371774 147922 371842 147978
rect 371898 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 402438 147978
rect 402494 147922 402562 147978
rect 402618 147922 433158 147978
rect 433214 147922 433282 147978
rect 433338 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 79878 136350
rect 79934 136294 80002 136350
rect 80058 136294 110598 136350
rect 110654 136294 110722 136350
rect 110778 136294 141318 136350
rect 141374 136294 141442 136350
rect 141498 136294 172038 136350
rect 172094 136294 172162 136350
rect 172218 136294 202758 136350
rect 202814 136294 202882 136350
rect 202938 136294 233478 136350
rect 233534 136294 233602 136350
rect 233658 136294 264198 136350
rect 264254 136294 264322 136350
rect 264378 136294 294918 136350
rect 294974 136294 295042 136350
rect 295098 136294 325638 136350
rect 325694 136294 325762 136350
rect 325818 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 356358 136350
rect 356414 136294 356482 136350
rect 356538 136294 366970 136350
rect 367026 136294 367094 136350
rect 367150 136294 367218 136350
rect 367274 136294 367342 136350
rect 367398 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 387078 136350
rect 387134 136294 387202 136350
rect 387258 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 417798 136350
rect 417854 136294 417922 136350
rect 417978 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 79878 136226
rect 79934 136170 80002 136226
rect 80058 136170 110598 136226
rect 110654 136170 110722 136226
rect 110778 136170 141318 136226
rect 141374 136170 141442 136226
rect 141498 136170 172038 136226
rect 172094 136170 172162 136226
rect 172218 136170 202758 136226
rect 202814 136170 202882 136226
rect 202938 136170 233478 136226
rect 233534 136170 233602 136226
rect 233658 136170 264198 136226
rect 264254 136170 264322 136226
rect 264378 136170 294918 136226
rect 294974 136170 295042 136226
rect 295098 136170 325638 136226
rect 325694 136170 325762 136226
rect 325818 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 356358 136226
rect 356414 136170 356482 136226
rect 356538 136170 366970 136226
rect 367026 136170 367094 136226
rect 367150 136170 367218 136226
rect 367274 136170 367342 136226
rect 367398 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 387078 136226
rect 387134 136170 387202 136226
rect 387258 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 417798 136226
rect 417854 136170 417922 136226
rect 417978 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 79878 136102
rect 79934 136046 80002 136102
rect 80058 136046 110598 136102
rect 110654 136046 110722 136102
rect 110778 136046 141318 136102
rect 141374 136046 141442 136102
rect 141498 136046 172038 136102
rect 172094 136046 172162 136102
rect 172218 136046 202758 136102
rect 202814 136046 202882 136102
rect 202938 136046 233478 136102
rect 233534 136046 233602 136102
rect 233658 136046 264198 136102
rect 264254 136046 264322 136102
rect 264378 136046 294918 136102
rect 294974 136046 295042 136102
rect 295098 136046 325638 136102
rect 325694 136046 325762 136102
rect 325818 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 356358 136102
rect 356414 136046 356482 136102
rect 356538 136046 366970 136102
rect 367026 136046 367094 136102
rect 367150 136046 367218 136102
rect 367274 136046 367342 136102
rect 367398 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 387078 136102
rect 387134 136046 387202 136102
rect 387258 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 417798 136102
rect 417854 136046 417922 136102
rect 417978 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 79878 135978
rect 79934 135922 80002 135978
rect 80058 135922 110598 135978
rect 110654 135922 110722 135978
rect 110778 135922 141318 135978
rect 141374 135922 141442 135978
rect 141498 135922 172038 135978
rect 172094 135922 172162 135978
rect 172218 135922 202758 135978
rect 202814 135922 202882 135978
rect 202938 135922 233478 135978
rect 233534 135922 233602 135978
rect 233658 135922 264198 135978
rect 264254 135922 264322 135978
rect 264378 135922 294918 135978
rect 294974 135922 295042 135978
rect 295098 135922 325638 135978
rect 325694 135922 325762 135978
rect 325818 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 356358 135978
rect 356414 135922 356482 135978
rect 356538 135922 366970 135978
rect 367026 135922 367094 135978
rect 367150 135922 367218 135978
rect 367274 135922 367342 135978
rect 367398 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 387078 135978
rect 387134 135922 387202 135978
rect 387258 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 417798 135978
rect 417854 135922 417922 135978
rect 417978 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 64518 130350
rect 64574 130294 64642 130350
rect 64698 130294 95238 130350
rect 95294 130294 95362 130350
rect 95418 130294 125958 130350
rect 126014 130294 126082 130350
rect 126138 130294 156678 130350
rect 156734 130294 156802 130350
rect 156858 130294 187398 130350
rect 187454 130294 187522 130350
rect 187578 130294 218118 130350
rect 218174 130294 218242 130350
rect 218298 130294 248838 130350
rect 248894 130294 248962 130350
rect 249018 130294 279558 130350
rect 279614 130294 279682 130350
rect 279738 130294 310278 130350
rect 310334 130294 310402 130350
rect 310458 130294 340998 130350
rect 341054 130294 341122 130350
rect 341178 130294 363250 130350
rect 363306 130294 363374 130350
rect 363430 130294 363498 130350
rect 363554 130294 363622 130350
rect 363678 130294 371718 130350
rect 371774 130294 371842 130350
rect 371898 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 402438 130350
rect 402494 130294 402562 130350
rect 402618 130294 433158 130350
rect 433214 130294 433282 130350
rect 433338 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 64518 130226
rect 64574 130170 64642 130226
rect 64698 130170 95238 130226
rect 95294 130170 95362 130226
rect 95418 130170 125958 130226
rect 126014 130170 126082 130226
rect 126138 130170 156678 130226
rect 156734 130170 156802 130226
rect 156858 130170 187398 130226
rect 187454 130170 187522 130226
rect 187578 130170 218118 130226
rect 218174 130170 218242 130226
rect 218298 130170 248838 130226
rect 248894 130170 248962 130226
rect 249018 130170 279558 130226
rect 279614 130170 279682 130226
rect 279738 130170 310278 130226
rect 310334 130170 310402 130226
rect 310458 130170 340998 130226
rect 341054 130170 341122 130226
rect 341178 130170 363250 130226
rect 363306 130170 363374 130226
rect 363430 130170 363498 130226
rect 363554 130170 363622 130226
rect 363678 130170 371718 130226
rect 371774 130170 371842 130226
rect 371898 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 402438 130226
rect 402494 130170 402562 130226
rect 402618 130170 433158 130226
rect 433214 130170 433282 130226
rect 433338 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 64518 130102
rect 64574 130046 64642 130102
rect 64698 130046 95238 130102
rect 95294 130046 95362 130102
rect 95418 130046 125958 130102
rect 126014 130046 126082 130102
rect 126138 130046 156678 130102
rect 156734 130046 156802 130102
rect 156858 130046 187398 130102
rect 187454 130046 187522 130102
rect 187578 130046 218118 130102
rect 218174 130046 218242 130102
rect 218298 130046 248838 130102
rect 248894 130046 248962 130102
rect 249018 130046 279558 130102
rect 279614 130046 279682 130102
rect 279738 130046 310278 130102
rect 310334 130046 310402 130102
rect 310458 130046 340998 130102
rect 341054 130046 341122 130102
rect 341178 130046 363250 130102
rect 363306 130046 363374 130102
rect 363430 130046 363498 130102
rect 363554 130046 363622 130102
rect 363678 130046 371718 130102
rect 371774 130046 371842 130102
rect 371898 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 402438 130102
rect 402494 130046 402562 130102
rect 402618 130046 433158 130102
rect 433214 130046 433282 130102
rect 433338 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 64518 129978
rect 64574 129922 64642 129978
rect 64698 129922 95238 129978
rect 95294 129922 95362 129978
rect 95418 129922 125958 129978
rect 126014 129922 126082 129978
rect 126138 129922 156678 129978
rect 156734 129922 156802 129978
rect 156858 129922 187398 129978
rect 187454 129922 187522 129978
rect 187578 129922 218118 129978
rect 218174 129922 218242 129978
rect 218298 129922 248838 129978
rect 248894 129922 248962 129978
rect 249018 129922 279558 129978
rect 279614 129922 279682 129978
rect 279738 129922 310278 129978
rect 310334 129922 310402 129978
rect 310458 129922 340998 129978
rect 341054 129922 341122 129978
rect 341178 129922 363250 129978
rect 363306 129922 363374 129978
rect 363430 129922 363498 129978
rect 363554 129922 363622 129978
rect 363678 129922 371718 129978
rect 371774 129922 371842 129978
rect 371898 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 402438 129978
rect 402494 129922 402562 129978
rect 402618 129922 433158 129978
rect 433214 129922 433282 129978
rect 433338 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 79878 118350
rect 79934 118294 80002 118350
rect 80058 118294 110598 118350
rect 110654 118294 110722 118350
rect 110778 118294 141318 118350
rect 141374 118294 141442 118350
rect 141498 118294 172038 118350
rect 172094 118294 172162 118350
rect 172218 118294 202758 118350
rect 202814 118294 202882 118350
rect 202938 118294 233478 118350
rect 233534 118294 233602 118350
rect 233658 118294 264198 118350
rect 264254 118294 264322 118350
rect 264378 118294 294918 118350
rect 294974 118294 295042 118350
rect 295098 118294 325638 118350
rect 325694 118294 325762 118350
rect 325818 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 356358 118350
rect 356414 118294 356482 118350
rect 356538 118294 366970 118350
rect 367026 118294 367094 118350
rect 367150 118294 367218 118350
rect 367274 118294 367342 118350
rect 367398 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 387078 118350
rect 387134 118294 387202 118350
rect 387258 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 417798 118350
rect 417854 118294 417922 118350
rect 417978 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 79878 118226
rect 79934 118170 80002 118226
rect 80058 118170 110598 118226
rect 110654 118170 110722 118226
rect 110778 118170 141318 118226
rect 141374 118170 141442 118226
rect 141498 118170 172038 118226
rect 172094 118170 172162 118226
rect 172218 118170 202758 118226
rect 202814 118170 202882 118226
rect 202938 118170 233478 118226
rect 233534 118170 233602 118226
rect 233658 118170 264198 118226
rect 264254 118170 264322 118226
rect 264378 118170 294918 118226
rect 294974 118170 295042 118226
rect 295098 118170 325638 118226
rect 325694 118170 325762 118226
rect 325818 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 356358 118226
rect 356414 118170 356482 118226
rect 356538 118170 366970 118226
rect 367026 118170 367094 118226
rect 367150 118170 367218 118226
rect 367274 118170 367342 118226
rect 367398 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 387078 118226
rect 387134 118170 387202 118226
rect 387258 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 417798 118226
rect 417854 118170 417922 118226
rect 417978 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 79878 118102
rect 79934 118046 80002 118102
rect 80058 118046 110598 118102
rect 110654 118046 110722 118102
rect 110778 118046 141318 118102
rect 141374 118046 141442 118102
rect 141498 118046 172038 118102
rect 172094 118046 172162 118102
rect 172218 118046 202758 118102
rect 202814 118046 202882 118102
rect 202938 118046 233478 118102
rect 233534 118046 233602 118102
rect 233658 118046 264198 118102
rect 264254 118046 264322 118102
rect 264378 118046 294918 118102
rect 294974 118046 295042 118102
rect 295098 118046 325638 118102
rect 325694 118046 325762 118102
rect 325818 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 356358 118102
rect 356414 118046 356482 118102
rect 356538 118046 366970 118102
rect 367026 118046 367094 118102
rect 367150 118046 367218 118102
rect 367274 118046 367342 118102
rect 367398 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 387078 118102
rect 387134 118046 387202 118102
rect 387258 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 417798 118102
rect 417854 118046 417922 118102
rect 417978 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 79878 117978
rect 79934 117922 80002 117978
rect 80058 117922 110598 117978
rect 110654 117922 110722 117978
rect 110778 117922 141318 117978
rect 141374 117922 141442 117978
rect 141498 117922 172038 117978
rect 172094 117922 172162 117978
rect 172218 117922 202758 117978
rect 202814 117922 202882 117978
rect 202938 117922 233478 117978
rect 233534 117922 233602 117978
rect 233658 117922 264198 117978
rect 264254 117922 264322 117978
rect 264378 117922 294918 117978
rect 294974 117922 295042 117978
rect 295098 117922 325638 117978
rect 325694 117922 325762 117978
rect 325818 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 356358 117978
rect 356414 117922 356482 117978
rect 356538 117922 366970 117978
rect 367026 117922 367094 117978
rect 367150 117922 367218 117978
rect 367274 117922 367342 117978
rect 367398 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 387078 117978
rect 387134 117922 387202 117978
rect 387258 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 417798 117978
rect 417854 117922 417922 117978
rect 417978 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 64518 112350
rect 64574 112294 64642 112350
rect 64698 112294 95238 112350
rect 95294 112294 95362 112350
rect 95418 112294 125958 112350
rect 126014 112294 126082 112350
rect 126138 112294 156678 112350
rect 156734 112294 156802 112350
rect 156858 112294 187398 112350
rect 187454 112294 187522 112350
rect 187578 112294 218118 112350
rect 218174 112294 218242 112350
rect 218298 112294 248838 112350
rect 248894 112294 248962 112350
rect 249018 112294 279558 112350
rect 279614 112294 279682 112350
rect 279738 112294 310278 112350
rect 310334 112294 310402 112350
rect 310458 112294 340998 112350
rect 341054 112294 341122 112350
rect 341178 112294 363250 112350
rect 363306 112294 363374 112350
rect 363430 112294 363498 112350
rect 363554 112294 363622 112350
rect 363678 112294 371718 112350
rect 371774 112294 371842 112350
rect 371898 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 402438 112350
rect 402494 112294 402562 112350
rect 402618 112294 433158 112350
rect 433214 112294 433282 112350
rect 433338 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 64518 112226
rect 64574 112170 64642 112226
rect 64698 112170 95238 112226
rect 95294 112170 95362 112226
rect 95418 112170 125958 112226
rect 126014 112170 126082 112226
rect 126138 112170 156678 112226
rect 156734 112170 156802 112226
rect 156858 112170 187398 112226
rect 187454 112170 187522 112226
rect 187578 112170 218118 112226
rect 218174 112170 218242 112226
rect 218298 112170 248838 112226
rect 248894 112170 248962 112226
rect 249018 112170 279558 112226
rect 279614 112170 279682 112226
rect 279738 112170 310278 112226
rect 310334 112170 310402 112226
rect 310458 112170 340998 112226
rect 341054 112170 341122 112226
rect 341178 112170 363250 112226
rect 363306 112170 363374 112226
rect 363430 112170 363498 112226
rect 363554 112170 363622 112226
rect 363678 112170 371718 112226
rect 371774 112170 371842 112226
rect 371898 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 402438 112226
rect 402494 112170 402562 112226
rect 402618 112170 433158 112226
rect 433214 112170 433282 112226
rect 433338 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 64518 112102
rect 64574 112046 64642 112102
rect 64698 112046 95238 112102
rect 95294 112046 95362 112102
rect 95418 112046 125958 112102
rect 126014 112046 126082 112102
rect 126138 112046 156678 112102
rect 156734 112046 156802 112102
rect 156858 112046 187398 112102
rect 187454 112046 187522 112102
rect 187578 112046 218118 112102
rect 218174 112046 218242 112102
rect 218298 112046 248838 112102
rect 248894 112046 248962 112102
rect 249018 112046 279558 112102
rect 279614 112046 279682 112102
rect 279738 112046 310278 112102
rect 310334 112046 310402 112102
rect 310458 112046 340998 112102
rect 341054 112046 341122 112102
rect 341178 112046 363250 112102
rect 363306 112046 363374 112102
rect 363430 112046 363498 112102
rect 363554 112046 363622 112102
rect 363678 112046 371718 112102
rect 371774 112046 371842 112102
rect 371898 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 402438 112102
rect 402494 112046 402562 112102
rect 402618 112046 433158 112102
rect 433214 112046 433282 112102
rect 433338 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 64518 111978
rect 64574 111922 64642 111978
rect 64698 111922 95238 111978
rect 95294 111922 95362 111978
rect 95418 111922 125958 111978
rect 126014 111922 126082 111978
rect 126138 111922 156678 111978
rect 156734 111922 156802 111978
rect 156858 111922 187398 111978
rect 187454 111922 187522 111978
rect 187578 111922 218118 111978
rect 218174 111922 218242 111978
rect 218298 111922 248838 111978
rect 248894 111922 248962 111978
rect 249018 111922 279558 111978
rect 279614 111922 279682 111978
rect 279738 111922 310278 111978
rect 310334 111922 310402 111978
rect 310458 111922 340998 111978
rect 341054 111922 341122 111978
rect 341178 111922 363250 111978
rect 363306 111922 363374 111978
rect 363430 111922 363498 111978
rect 363554 111922 363622 111978
rect 363678 111922 371718 111978
rect 371774 111922 371842 111978
rect 371898 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 402438 111978
rect 402494 111922 402562 111978
rect 402618 111922 433158 111978
rect 433214 111922 433282 111978
rect 433338 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 79878 100350
rect 79934 100294 80002 100350
rect 80058 100294 110598 100350
rect 110654 100294 110722 100350
rect 110778 100294 141318 100350
rect 141374 100294 141442 100350
rect 141498 100294 172038 100350
rect 172094 100294 172162 100350
rect 172218 100294 202758 100350
rect 202814 100294 202882 100350
rect 202938 100294 233478 100350
rect 233534 100294 233602 100350
rect 233658 100294 264198 100350
rect 264254 100294 264322 100350
rect 264378 100294 294918 100350
rect 294974 100294 295042 100350
rect 295098 100294 325638 100350
rect 325694 100294 325762 100350
rect 325818 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 356358 100350
rect 356414 100294 356482 100350
rect 356538 100294 366970 100350
rect 367026 100294 367094 100350
rect 367150 100294 367218 100350
rect 367274 100294 367342 100350
rect 367398 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 387078 100350
rect 387134 100294 387202 100350
rect 387258 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 417798 100350
rect 417854 100294 417922 100350
rect 417978 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 79878 100226
rect 79934 100170 80002 100226
rect 80058 100170 110598 100226
rect 110654 100170 110722 100226
rect 110778 100170 141318 100226
rect 141374 100170 141442 100226
rect 141498 100170 172038 100226
rect 172094 100170 172162 100226
rect 172218 100170 202758 100226
rect 202814 100170 202882 100226
rect 202938 100170 233478 100226
rect 233534 100170 233602 100226
rect 233658 100170 264198 100226
rect 264254 100170 264322 100226
rect 264378 100170 294918 100226
rect 294974 100170 295042 100226
rect 295098 100170 325638 100226
rect 325694 100170 325762 100226
rect 325818 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 356358 100226
rect 356414 100170 356482 100226
rect 356538 100170 366970 100226
rect 367026 100170 367094 100226
rect 367150 100170 367218 100226
rect 367274 100170 367342 100226
rect 367398 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 387078 100226
rect 387134 100170 387202 100226
rect 387258 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 417798 100226
rect 417854 100170 417922 100226
rect 417978 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 79878 100102
rect 79934 100046 80002 100102
rect 80058 100046 110598 100102
rect 110654 100046 110722 100102
rect 110778 100046 141318 100102
rect 141374 100046 141442 100102
rect 141498 100046 172038 100102
rect 172094 100046 172162 100102
rect 172218 100046 202758 100102
rect 202814 100046 202882 100102
rect 202938 100046 233478 100102
rect 233534 100046 233602 100102
rect 233658 100046 264198 100102
rect 264254 100046 264322 100102
rect 264378 100046 294918 100102
rect 294974 100046 295042 100102
rect 295098 100046 325638 100102
rect 325694 100046 325762 100102
rect 325818 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 356358 100102
rect 356414 100046 356482 100102
rect 356538 100046 366970 100102
rect 367026 100046 367094 100102
rect 367150 100046 367218 100102
rect 367274 100046 367342 100102
rect 367398 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 387078 100102
rect 387134 100046 387202 100102
rect 387258 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 417798 100102
rect 417854 100046 417922 100102
rect 417978 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 79878 99978
rect 79934 99922 80002 99978
rect 80058 99922 110598 99978
rect 110654 99922 110722 99978
rect 110778 99922 141318 99978
rect 141374 99922 141442 99978
rect 141498 99922 172038 99978
rect 172094 99922 172162 99978
rect 172218 99922 202758 99978
rect 202814 99922 202882 99978
rect 202938 99922 233478 99978
rect 233534 99922 233602 99978
rect 233658 99922 264198 99978
rect 264254 99922 264322 99978
rect 264378 99922 294918 99978
rect 294974 99922 295042 99978
rect 295098 99922 325638 99978
rect 325694 99922 325762 99978
rect 325818 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 356358 99978
rect 356414 99922 356482 99978
rect 356538 99922 366970 99978
rect 367026 99922 367094 99978
rect 367150 99922 367218 99978
rect 367274 99922 367342 99978
rect 367398 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 387078 99978
rect 387134 99922 387202 99978
rect 387258 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 417798 99978
rect 417854 99922 417922 99978
rect 417978 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 64518 94350
rect 64574 94294 64642 94350
rect 64698 94294 95238 94350
rect 95294 94294 95362 94350
rect 95418 94294 125958 94350
rect 126014 94294 126082 94350
rect 126138 94294 156678 94350
rect 156734 94294 156802 94350
rect 156858 94294 187398 94350
rect 187454 94294 187522 94350
rect 187578 94294 218118 94350
rect 218174 94294 218242 94350
rect 218298 94294 248838 94350
rect 248894 94294 248962 94350
rect 249018 94294 279558 94350
rect 279614 94294 279682 94350
rect 279738 94294 310278 94350
rect 310334 94294 310402 94350
rect 310458 94294 340998 94350
rect 341054 94294 341122 94350
rect 341178 94294 363250 94350
rect 363306 94294 363374 94350
rect 363430 94294 363498 94350
rect 363554 94294 363622 94350
rect 363678 94294 371718 94350
rect 371774 94294 371842 94350
rect 371898 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 402438 94350
rect 402494 94294 402562 94350
rect 402618 94294 433158 94350
rect 433214 94294 433282 94350
rect 433338 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 64518 94226
rect 64574 94170 64642 94226
rect 64698 94170 95238 94226
rect 95294 94170 95362 94226
rect 95418 94170 125958 94226
rect 126014 94170 126082 94226
rect 126138 94170 156678 94226
rect 156734 94170 156802 94226
rect 156858 94170 187398 94226
rect 187454 94170 187522 94226
rect 187578 94170 218118 94226
rect 218174 94170 218242 94226
rect 218298 94170 248838 94226
rect 248894 94170 248962 94226
rect 249018 94170 279558 94226
rect 279614 94170 279682 94226
rect 279738 94170 310278 94226
rect 310334 94170 310402 94226
rect 310458 94170 340998 94226
rect 341054 94170 341122 94226
rect 341178 94170 363250 94226
rect 363306 94170 363374 94226
rect 363430 94170 363498 94226
rect 363554 94170 363622 94226
rect 363678 94170 371718 94226
rect 371774 94170 371842 94226
rect 371898 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 402438 94226
rect 402494 94170 402562 94226
rect 402618 94170 433158 94226
rect 433214 94170 433282 94226
rect 433338 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 64518 94102
rect 64574 94046 64642 94102
rect 64698 94046 95238 94102
rect 95294 94046 95362 94102
rect 95418 94046 125958 94102
rect 126014 94046 126082 94102
rect 126138 94046 156678 94102
rect 156734 94046 156802 94102
rect 156858 94046 187398 94102
rect 187454 94046 187522 94102
rect 187578 94046 218118 94102
rect 218174 94046 218242 94102
rect 218298 94046 248838 94102
rect 248894 94046 248962 94102
rect 249018 94046 279558 94102
rect 279614 94046 279682 94102
rect 279738 94046 310278 94102
rect 310334 94046 310402 94102
rect 310458 94046 340998 94102
rect 341054 94046 341122 94102
rect 341178 94046 363250 94102
rect 363306 94046 363374 94102
rect 363430 94046 363498 94102
rect 363554 94046 363622 94102
rect 363678 94046 371718 94102
rect 371774 94046 371842 94102
rect 371898 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 402438 94102
rect 402494 94046 402562 94102
rect 402618 94046 433158 94102
rect 433214 94046 433282 94102
rect 433338 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 64518 93978
rect 64574 93922 64642 93978
rect 64698 93922 95238 93978
rect 95294 93922 95362 93978
rect 95418 93922 125958 93978
rect 126014 93922 126082 93978
rect 126138 93922 156678 93978
rect 156734 93922 156802 93978
rect 156858 93922 187398 93978
rect 187454 93922 187522 93978
rect 187578 93922 218118 93978
rect 218174 93922 218242 93978
rect 218298 93922 248838 93978
rect 248894 93922 248962 93978
rect 249018 93922 279558 93978
rect 279614 93922 279682 93978
rect 279738 93922 310278 93978
rect 310334 93922 310402 93978
rect 310458 93922 340998 93978
rect 341054 93922 341122 93978
rect 341178 93922 363250 93978
rect 363306 93922 363374 93978
rect 363430 93922 363498 93978
rect 363554 93922 363622 93978
rect 363678 93922 371718 93978
rect 371774 93922 371842 93978
rect 371898 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 402438 93978
rect 402494 93922 402562 93978
rect 402618 93922 433158 93978
rect 433214 93922 433282 93978
rect 433338 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 79878 82350
rect 79934 82294 80002 82350
rect 80058 82294 110598 82350
rect 110654 82294 110722 82350
rect 110778 82294 141318 82350
rect 141374 82294 141442 82350
rect 141498 82294 172038 82350
rect 172094 82294 172162 82350
rect 172218 82294 202758 82350
rect 202814 82294 202882 82350
rect 202938 82294 233478 82350
rect 233534 82294 233602 82350
rect 233658 82294 264198 82350
rect 264254 82294 264322 82350
rect 264378 82294 294918 82350
rect 294974 82294 295042 82350
rect 295098 82294 325638 82350
rect 325694 82294 325762 82350
rect 325818 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 356358 82350
rect 356414 82294 356482 82350
rect 356538 82294 366970 82350
rect 367026 82294 367094 82350
rect 367150 82294 367218 82350
rect 367274 82294 367342 82350
rect 367398 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 387078 82350
rect 387134 82294 387202 82350
rect 387258 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 417798 82350
rect 417854 82294 417922 82350
rect 417978 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 79878 82226
rect 79934 82170 80002 82226
rect 80058 82170 110598 82226
rect 110654 82170 110722 82226
rect 110778 82170 141318 82226
rect 141374 82170 141442 82226
rect 141498 82170 172038 82226
rect 172094 82170 172162 82226
rect 172218 82170 202758 82226
rect 202814 82170 202882 82226
rect 202938 82170 233478 82226
rect 233534 82170 233602 82226
rect 233658 82170 264198 82226
rect 264254 82170 264322 82226
rect 264378 82170 294918 82226
rect 294974 82170 295042 82226
rect 295098 82170 325638 82226
rect 325694 82170 325762 82226
rect 325818 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 356358 82226
rect 356414 82170 356482 82226
rect 356538 82170 366970 82226
rect 367026 82170 367094 82226
rect 367150 82170 367218 82226
rect 367274 82170 367342 82226
rect 367398 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 387078 82226
rect 387134 82170 387202 82226
rect 387258 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 417798 82226
rect 417854 82170 417922 82226
rect 417978 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 79878 82102
rect 79934 82046 80002 82102
rect 80058 82046 110598 82102
rect 110654 82046 110722 82102
rect 110778 82046 141318 82102
rect 141374 82046 141442 82102
rect 141498 82046 172038 82102
rect 172094 82046 172162 82102
rect 172218 82046 202758 82102
rect 202814 82046 202882 82102
rect 202938 82046 233478 82102
rect 233534 82046 233602 82102
rect 233658 82046 264198 82102
rect 264254 82046 264322 82102
rect 264378 82046 294918 82102
rect 294974 82046 295042 82102
rect 295098 82046 325638 82102
rect 325694 82046 325762 82102
rect 325818 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 356358 82102
rect 356414 82046 356482 82102
rect 356538 82046 366970 82102
rect 367026 82046 367094 82102
rect 367150 82046 367218 82102
rect 367274 82046 367342 82102
rect 367398 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 387078 82102
rect 387134 82046 387202 82102
rect 387258 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 417798 82102
rect 417854 82046 417922 82102
rect 417978 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 79878 81978
rect 79934 81922 80002 81978
rect 80058 81922 110598 81978
rect 110654 81922 110722 81978
rect 110778 81922 141318 81978
rect 141374 81922 141442 81978
rect 141498 81922 172038 81978
rect 172094 81922 172162 81978
rect 172218 81922 202758 81978
rect 202814 81922 202882 81978
rect 202938 81922 233478 81978
rect 233534 81922 233602 81978
rect 233658 81922 264198 81978
rect 264254 81922 264322 81978
rect 264378 81922 294918 81978
rect 294974 81922 295042 81978
rect 295098 81922 325638 81978
rect 325694 81922 325762 81978
rect 325818 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 356358 81978
rect 356414 81922 356482 81978
rect 356538 81922 366970 81978
rect 367026 81922 367094 81978
rect 367150 81922 367218 81978
rect 367274 81922 367342 81978
rect 367398 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 387078 81978
rect 387134 81922 387202 81978
rect 387258 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 417798 81978
rect 417854 81922 417922 81978
rect 417978 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 64518 76350
rect 64574 76294 64642 76350
rect 64698 76294 95238 76350
rect 95294 76294 95362 76350
rect 95418 76294 125958 76350
rect 126014 76294 126082 76350
rect 126138 76294 156678 76350
rect 156734 76294 156802 76350
rect 156858 76294 187398 76350
rect 187454 76294 187522 76350
rect 187578 76294 218118 76350
rect 218174 76294 218242 76350
rect 218298 76294 248838 76350
rect 248894 76294 248962 76350
rect 249018 76294 279558 76350
rect 279614 76294 279682 76350
rect 279738 76294 310278 76350
rect 310334 76294 310402 76350
rect 310458 76294 340998 76350
rect 341054 76294 341122 76350
rect 341178 76294 363250 76350
rect 363306 76294 363374 76350
rect 363430 76294 363498 76350
rect 363554 76294 363622 76350
rect 363678 76294 371718 76350
rect 371774 76294 371842 76350
rect 371898 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 402438 76350
rect 402494 76294 402562 76350
rect 402618 76294 433158 76350
rect 433214 76294 433282 76350
rect 433338 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 64518 76226
rect 64574 76170 64642 76226
rect 64698 76170 95238 76226
rect 95294 76170 95362 76226
rect 95418 76170 125958 76226
rect 126014 76170 126082 76226
rect 126138 76170 156678 76226
rect 156734 76170 156802 76226
rect 156858 76170 187398 76226
rect 187454 76170 187522 76226
rect 187578 76170 218118 76226
rect 218174 76170 218242 76226
rect 218298 76170 248838 76226
rect 248894 76170 248962 76226
rect 249018 76170 279558 76226
rect 279614 76170 279682 76226
rect 279738 76170 310278 76226
rect 310334 76170 310402 76226
rect 310458 76170 340998 76226
rect 341054 76170 341122 76226
rect 341178 76170 363250 76226
rect 363306 76170 363374 76226
rect 363430 76170 363498 76226
rect 363554 76170 363622 76226
rect 363678 76170 371718 76226
rect 371774 76170 371842 76226
rect 371898 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 402438 76226
rect 402494 76170 402562 76226
rect 402618 76170 433158 76226
rect 433214 76170 433282 76226
rect 433338 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 64518 76102
rect 64574 76046 64642 76102
rect 64698 76046 95238 76102
rect 95294 76046 95362 76102
rect 95418 76046 125958 76102
rect 126014 76046 126082 76102
rect 126138 76046 156678 76102
rect 156734 76046 156802 76102
rect 156858 76046 187398 76102
rect 187454 76046 187522 76102
rect 187578 76046 218118 76102
rect 218174 76046 218242 76102
rect 218298 76046 248838 76102
rect 248894 76046 248962 76102
rect 249018 76046 279558 76102
rect 279614 76046 279682 76102
rect 279738 76046 310278 76102
rect 310334 76046 310402 76102
rect 310458 76046 340998 76102
rect 341054 76046 341122 76102
rect 341178 76046 363250 76102
rect 363306 76046 363374 76102
rect 363430 76046 363498 76102
rect 363554 76046 363622 76102
rect 363678 76046 371718 76102
rect 371774 76046 371842 76102
rect 371898 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 402438 76102
rect 402494 76046 402562 76102
rect 402618 76046 433158 76102
rect 433214 76046 433282 76102
rect 433338 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 64518 75978
rect 64574 75922 64642 75978
rect 64698 75922 95238 75978
rect 95294 75922 95362 75978
rect 95418 75922 125958 75978
rect 126014 75922 126082 75978
rect 126138 75922 156678 75978
rect 156734 75922 156802 75978
rect 156858 75922 187398 75978
rect 187454 75922 187522 75978
rect 187578 75922 218118 75978
rect 218174 75922 218242 75978
rect 218298 75922 248838 75978
rect 248894 75922 248962 75978
rect 249018 75922 279558 75978
rect 279614 75922 279682 75978
rect 279738 75922 310278 75978
rect 310334 75922 310402 75978
rect 310458 75922 340998 75978
rect 341054 75922 341122 75978
rect 341178 75922 363250 75978
rect 363306 75922 363374 75978
rect 363430 75922 363498 75978
rect 363554 75922 363622 75978
rect 363678 75922 371718 75978
rect 371774 75922 371842 75978
rect 371898 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 402438 75978
rect 402494 75922 402562 75978
rect 402618 75922 433158 75978
rect 433214 75922 433282 75978
rect 433338 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 79878 64350
rect 79934 64294 80002 64350
rect 80058 64294 110598 64350
rect 110654 64294 110722 64350
rect 110778 64294 141318 64350
rect 141374 64294 141442 64350
rect 141498 64294 172038 64350
rect 172094 64294 172162 64350
rect 172218 64294 202758 64350
rect 202814 64294 202882 64350
rect 202938 64294 233478 64350
rect 233534 64294 233602 64350
rect 233658 64294 264198 64350
rect 264254 64294 264322 64350
rect 264378 64294 294918 64350
rect 294974 64294 295042 64350
rect 295098 64294 325638 64350
rect 325694 64294 325762 64350
rect 325818 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 356358 64350
rect 356414 64294 356482 64350
rect 356538 64294 366970 64350
rect 367026 64294 367094 64350
rect 367150 64294 367218 64350
rect 367274 64294 367342 64350
rect 367398 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 387078 64350
rect 387134 64294 387202 64350
rect 387258 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 417798 64350
rect 417854 64294 417922 64350
rect 417978 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 79878 64226
rect 79934 64170 80002 64226
rect 80058 64170 110598 64226
rect 110654 64170 110722 64226
rect 110778 64170 141318 64226
rect 141374 64170 141442 64226
rect 141498 64170 172038 64226
rect 172094 64170 172162 64226
rect 172218 64170 202758 64226
rect 202814 64170 202882 64226
rect 202938 64170 233478 64226
rect 233534 64170 233602 64226
rect 233658 64170 264198 64226
rect 264254 64170 264322 64226
rect 264378 64170 294918 64226
rect 294974 64170 295042 64226
rect 295098 64170 325638 64226
rect 325694 64170 325762 64226
rect 325818 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 356358 64226
rect 356414 64170 356482 64226
rect 356538 64170 366970 64226
rect 367026 64170 367094 64226
rect 367150 64170 367218 64226
rect 367274 64170 367342 64226
rect 367398 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 387078 64226
rect 387134 64170 387202 64226
rect 387258 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 417798 64226
rect 417854 64170 417922 64226
rect 417978 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 79878 64102
rect 79934 64046 80002 64102
rect 80058 64046 110598 64102
rect 110654 64046 110722 64102
rect 110778 64046 141318 64102
rect 141374 64046 141442 64102
rect 141498 64046 172038 64102
rect 172094 64046 172162 64102
rect 172218 64046 202758 64102
rect 202814 64046 202882 64102
rect 202938 64046 233478 64102
rect 233534 64046 233602 64102
rect 233658 64046 264198 64102
rect 264254 64046 264322 64102
rect 264378 64046 294918 64102
rect 294974 64046 295042 64102
rect 295098 64046 325638 64102
rect 325694 64046 325762 64102
rect 325818 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 356358 64102
rect 356414 64046 356482 64102
rect 356538 64046 366970 64102
rect 367026 64046 367094 64102
rect 367150 64046 367218 64102
rect 367274 64046 367342 64102
rect 367398 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 387078 64102
rect 387134 64046 387202 64102
rect 387258 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 417798 64102
rect 417854 64046 417922 64102
rect 417978 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 79878 63978
rect 79934 63922 80002 63978
rect 80058 63922 110598 63978
rect 110654 63922 110722 63978
rect 110778 63922 141318 63978
rect 141374 63922 141442 63978
rect 141498 63922 172038 63978
rect 172094 63922 172162 63978
rect 172218 63922 202758 63978
rect 202814 63922 202882 63978
rect 202938 63922 233478 63978
rect 233534 63922 233602 63978
rect 233658 63922 264198 63978
rect 264254 63922 264322 63978
rect 264378 63922 294918 63978
rect 294974 63922 295042 63978
rect 295098 63922 325638 63978
rect 325694 63922 325762 63978
rect 325818 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 356358 63978
rect 356414 63922 356482 63978
rect 356538 63922 366970 63978
rect 367026 63922 367094 63978
rect 367150 63922 367218 63978
rect 367274 63922 367342 63978
rect 367398 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 387078 63978
rect 387134 63922 387202 63978
rect 387258 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 417798 63978
rect 417854 63922 417922 63978
rect 417978 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 219250 58350
rect 219306 58294 219374 58350
rect 219430 58294 219498 58350
rect 219554 58294 219622 58350
rect 219678 58294 237250 58350
rect 237306 58294 237374 58350
rect 237430 58294 237498 58350
rect 237554 58294 237622 58350
rect 237678 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 363250 58350
rect 363306 58294 363374 58350
rect 363430 58294 363498 58350
rect 363554 58294 363622 58350
rect 363678 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 219250 58226
rect 219306 58170 219374 58226
rect 219430 58170 219498 58226
rect 219554 58170 219622 58226
rect 219678 58170 237250 58226
rect 237306 58170 237374 58226
rect 237430 58170 237498 58226
rect 237554 58170 237622 58226
rect 237678 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 363250 58226
rect 363306 58170 363374 58226
rect 363430 58170 363498 58226
rect 363554 58170 363622 58226
rect 363678 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 219250 58102
rect 219306 58046 219374 58102
rect 219430 58046 219498 58102
rect 219554 58046 219622 58102
rect 219678 58046 237250 58102
rect 237306 58046 237374 58102
rect 237430 58046 237498 58102
rect 237554 58046 237622 58102
rect 237678 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 363250 58102
rect 363306 58046 363374 58102
rect 363430 58046 363498 58102
rect 363554 58046 363622 58102
rect 363678 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 219250 57978
rect 219306 57922 219374 57978
rect 219430 57922 219498 57978
rect 219554 57922 219622 57978
rect 219678 57922 237250 57978
rect 237306 57922 237374 57978
rect 237430 57922 237498 57978
rect 237554 57922 237622 57978
rect 237678 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 363250 57978
rect 363306 57922 363374 57978
rect 363430 57922 363498 57978
rect 363554 57922 363622 57978
rect 363678 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 222970 46350
rect 223026 46294 223094 46350
rect 223150 46294 223218 46350
rect 223274 46294 223342 46350
rect 223398 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 366970 46350
rect 367026 46294 367094 46350
rect 367150 46294 367218 46350
rect 367274 46294 367342 46350
rect 367398 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 222970 46226
rect 223026 46170 223094 46226
rect 223150 46170 223218 46226
rect 223274 46170 223342 46226
rect 223398 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 366970 46226
rect 367026 46170 367094 46226
rect 367150 46170 367218 46226
rect 367274 46170 367342 46226
rect 367398 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 222970 46102
rect 223026 46046 223094 46102
rect 223150 46046 223218 46102
rect 223274 46046 223342 46102
rect 223398 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 366970 46102
rect 367026 46046 367094 46102
rect 367150 46046 367218 46102
rect 367274 46046 367342 46102
rect 367398 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 222970 45978
rect 223026 45922 223094 45978
rect 223150 45922 223218 45978
rect 223274 45922 223342 45978
rect 223398 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 366970 45978
rect 367026 45922 367094 45978
rect 367150 45922 367218 45978
rect 367274 45922 367342 45978
rect 367398 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 219250 40350
rect 219306 40294 219374 40350
rect 219430 40294 219498 40350
rect 219554 40294 219622 40350
rect 219678 40294 237250 40350
rect 237306 40294 237374 40350
rect 237430 40294 237498 40350
rect 237554 40294 237622 40350
rect 237678 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 219250 40226
rect 219306 40170 219374 40226
rect 219430 40170 219498 40226
rect 219554 40170 219622 40226
rect 219678 40170 237250 40226
rect 237306 40170 237374 40226
rect 237430 40170 237498 40226
rect 237554 40170 237622 40226
rect 237678 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 219250 40102
rect 219306 40046 219374 40102
rect 219430 40046 219498 40102
rect 219554 40046 219622 40102
rect 219678 40046 237250 40102
rect 237306 40046 237374 40102
rect 237430 40046 237498 40102
rect 237554 40046 237622 40102
rect 237678 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 219250 39978
rect 219306 39922 219374 39978
rect 219430 39922 219498 39978
rect 219554 39922 219622 39978
rect 219678 39922 237250 39978
rect 237306 39922 237374 39978
rect 237430 39922 237498 39978
rect 237554 39922 237622 39978
rect 237678 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use user_proj  mprj
timestamp 0
transform 1 0 60000 0 1 60000
box 1138 0 378560 380000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 436006 75774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 436006 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 436006 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 436006 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 436006 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 436006 165774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 436006 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 436006 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 436006 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 436006 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 436006 255774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 436006 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 436006 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 436006 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 436006 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 59082 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 436006 345774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 61020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 438436 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 436006 61494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 436006 79494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 436006 97494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 436006 115494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 436006 133494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 436006 151494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 436006 169494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 438436 187494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 436006 205494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 -1644 223494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 436006 223494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 -1644 241494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 436006 241494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 -1644 259494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 436006 259494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 -1644 277494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 436006 277494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 -1644 295494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 438436 295494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 -1644 313494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 436006 313494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 -1644 331494 59082 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 436006 331494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 -1644 349494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 -1644 367494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 435650 436322 435650 436322 0 vdd
rlabel via4 439370 424322 439370 424322 0 vss
rlabel metal3 594986 7336 594986 7336 0 io_in[0]
rlabel metal3 594370 403816 594370 403816 0 io_in[10]
rlabel metal2 173362 439880 173362 439880 0 io_in[11]
rlabel metal3 595672 482496 595672 482496 0 io_in[12]
rlabel metal3 594426 522536 594426 522536 0 io_in[13]
rlabel metal3 594370 562184 594370 562184 0 io_in[14]
rlabel metal2 212226 439880 212226 439880 0 io_in[15]
rlabel metal2 518504 594426 518504 594426 0 io_in[16]
rlabel metal2 451640 594552 451640 594552 0 io_in[17]
rlabel metal2 386120 593138 386120 593138 0 io_in[18]
rlabel metal3 284816 503160 284816 503160 0 io_in[19]
rlabel metal2 76216 442582 76216 442582 0 io_in[1]
rlabel metal2 260946 439880 260946 439880 0 io_in[20]
rlabel metal2 189000 531776 189000 531776 0 io_in[21]
rlabel metal2 121184 588000 121184 588000 0 io_in[22]
rlabel metal2 55384 594482 55384 594482 0 io_in[23]
rlabel metal3 392 586712 392 586712 0 io_in[24]
rlabel metal3 392 544544 392 544544 0 io_in[25]
rlabel metal3 11760 502432 11760 502432 0 io_in[26]
rlabel metal3 392 459424 392 459424 0 io_in[27]
rlabel metal3 392 417200 392 417200 0 io_in[28]
rlabel metal3 392 375032 392 375032 0 io_in[29]
rlabel metal3 594594 86632 594594 86632 0 io_in[2]
rlabel metal3 392 332864 392 332864 0 io_in[30]
rlabel metal3 3150 291032 3150 291032 0 io_in[31]
rlabel metal3 392 247688 392 247688 0 io_in[32]
rlabel metal3 392 205520 392 205520 0 io_in[33]
rlabel metal3 392 163352 392 163352 0 io_in[34]
rlabel metal3 4830 121688 4830 121688 0 io_in[35]
rlabel metal3 11760 79072 11760 79072 0 io_in[36]
rlabel metal3 2702 36904 2702 36904 0 io_in[37]
rlabel metal3 594650 126280 594650 126280 0 io_in[3]
rlabel metal3 594762 165928 594762 165928 0 io_in[4]
rlabel metal3 588000 205184 588000 205184 0 io_in[5]
rlabel metal3 594818 245224 594818 245224 0 io_in[6]
rlabel metal3 594874 284872 594874 284872 0 io_in[7]
rlabel metal2 144018 439880 144018 439880 0 io_in[8]
rlabel metal3 595672 363384 595672 363384 0 io_in[9]
rlabel metal3 594426 33768 594426 33768 0 io_oeb[0]
rlabel metal2 167160 441966 167160 441966 0 io_oeb[10]
rlabel metal3 595672 469168 595672 469168 0 io_oeb[11]
rlabel metal2 194040 476728 194040 476728 0 io_oeb[12]
rlabel metal3 595672 548296 595672 548296 0 io_oeb[13]
rlabel metal3 595672 588280 595672 588280 0 io_oeb[14]
rlabel metal2 215474 439880 215474 439880 0 io_oeb[15]
rlabel metal2 474376 593082 474376 593082 0 io_oeb[16]
rlabel metal2 235298 439880 235298 439880 0 io_oeb[17]
rlabel metal2 244706 439880 244706 439880 0 io_oeb[18]
rlabel metal2 275688 588000 275688 588000 0 io_oeb[19]
rlabel metal3 594538 73416 594538 73416 0 io_oeb[1]
rlabel metal2 264194 439880 264194 439880 0 io_oeb[20]
rlabel metal2 143080 595672 143080 595672 0 io_oeb[21]
rlabel metal2 77336 519330 77336 519330 0 io_oeb[22]
rlabel metal2 10528 595672 10528 595672 0 io_oeb[23]
rlabel metal3 392 558320 392 558320 0 io_oeb[24]
rlabel metal3 2310 516600 2310 516600 0 io_oeb[25]
rlabel metal3 392 473984 392 473984 0 io_oeb[26]
rlabel metal3 11760 431872 11760 431872 0 io_oeb[27]
rlabel metal3 392 388808 392 388808 0 io_oeb[28]
rlabel metal3 392 346640 392 346640 0 io_oeb[29]
rlabel metal2 456120 279048 456120 279048 0 io_oeb[2]
rlabel metal3 392 304472 392 304472 0 io_oeb[30]
rlabel metal3 392 262304 392 262304 0 io_oeb[31]
rlabel metal3 5670 220472 5670 220472 0 io_oeb[32]
rlabel metal3 392 177128 392 177128 0 io_oeb[33]
rlabel metal3 392 134960 392 134960 0 io_oeb[34]
rlabel metal3 392 92792 392 92792 0 io_oeb[35]
rlabel metal3 392 50624 392 50624 0 io_oeb[36]
rlabel metal3 11760 8512 11760 8512 0 io_oeb[37]
rlabel metal3 594706 152712 594706 152712 0 io_oeb[3]
rlabel metal3 593082 192360 593082 192360 0 io_oeb[4]
rlabel metal2 118034 439880 118034 439880 0 io_oeb[5]
rlabel metal2 127946 439880 127946 439880 0 io_oeb[6]
rlabel metal3 588000 310968 588000 310968 0 io_oeb[7]
rlabel metal2 146216 448812 146216 448812 0 io_oeb[8]
rlabel metal3 595672 390040 595672 390040 0 io_oeb[9]
rlabel metal2 72968 440902 72968 440902 0 io_out[0]
rlabel metal2 170408 440958 170408 440958 0 io_out[10]
rlabel metal3 595672 455840 595672 455840 0 io_out[11]
rlabel metal3 595672 495824 595672 495824 0 io_out[12]
rlabel metal2 199234 439880 199234 439880 0 io_out[13]
rlabel metal3 595672 574952 595672 574952 0 io_out[14]
rlabel metal2 219128 441294 219128 441294 0 io_out[15]
rlabel metal2 495992 595672 495992 595672 0 io_out[16]
rlabel metal3 428904 590856 428904 590856 0 io_out[17]
rlabel metal2 364056 593082 364056 593082 0 io_out[18]
rlabel metal2 297584 595672 297584 595672 0 io_out[19]
rlabel metal2 496440 252952 496440 252952 0 io_out[1]
rlabel metal2 267498 439880 267498 439880 0 io_out[20]
rlabel metal2 165032 595672 165032 595672 0 io_out[21]
rlabel metal3 102256 591304 102256 591304 0 io_out[22]
rlabel metal2 33320 593082 33320 593082 0 io_out[23]
rlabel metal3 11760 572992 11760 572992 0 io_out[24]
rlabel metal3 3150 530712 3150 530712 0 io_out[25]
rlabel metal3 392 487760 392 487760 0 io_out[26]
rlabel metal3 392 445648 392 445648 0 io_out[27]
rlabel metal3 392 403424 392 403424 0 io_out[28]
rlabel metal3 11760 361312 11760 361312 0 io_out[29]
rlabel metal3 595672 99344 595672 99344 0 io_out[2]
rlabel metal3 392 318248 392 318248 0 io_out[30]
rlabel metal3 392 276080 392 276080 0 io_out[31]
rlabel metal3 392 233912 392 233912 0 io_out[32]
rlabel metal3 392 191744 392 191744 0 io_out[33]
rlabel metal3 11760 149632 11760 149632 0 io_out[34]
rlabel metal3 1470 107464 1470 107464 0 io_out[35]
rlabel metal3 392 64400 392 64400 0 io_out[36]
rlabel metal3 392 22232 392 22232 0 io_out[37]
rlabel metal2 100856 450324 100856 450324 0 io_out[3]
rlabel metal2 454440 310016 454440 310016 0 io_out[4]
rlabel metal3 588000 218512 588000 218512 0 io_out[5]
rlabel metal2 479640 352184 479640 352184 0 io_out[6]
rlabel metal2 141176 447622 141176 447622 0 io_out[7]
rlabel metal3 595672 336728 595672 336728 0 io_out[8]
rlabel metal3 595672 376712 595672 376712 0 io_out[9]
rlabel metal2 213192 3206 213192 3206 0 la_data_in[0]
rlabel metal2 269584 392 269584 392 0 la_data_in[10]
rlabel metal2 235914 60088 235914 60088 0 la_data_in[11]
rlabel metal3 239064 59416 239064 59416 0 la_data_in[12]
rlabel metal2 287448 4046 287448 4046 0 la_data_in[13]
rlabel metal2 293160 5782 293160 5782 0 la_data_in[14]
rlabel metal2 298088 392 298088 392 0 la_data_in[15]
rlabel metal2 286440 32144 286440 32144 0 la_data_in[16]
rlabel metal3 309288 4984 309288 4984 0 la_data_in[17]
rlabel metal2 315952 11760 315952 11760 0 la_data_in[18]
rlabel metal2 265762 60088 265762 60088 0 la_data_in[19]
rlabel metal2 218344 7952 218344 7952 0 la_data_in[1]
rlabel metal2 269290 60088 269290 60088 0 la_data_in[20]
rlabel metal2 332920 392 332920 392 0 la_data_in[21]
rlabel metal3 337008 5768 337008 5768 0 la_data_in[22]
rlabel metal2 344568 3206 344568 3206 0 la_data_in[23]
rlabel metal2 284242 60088 284242 60088 0 la_data_in[24]
rlabel metal2 355992 5670 355992 5670 0 la_data_in[25]
rlabel metal3 359352 8120 359352 8120 0 la_data_in[26]
rlabel metal2 362040 31360 362040 31360 0 la_data_in[27]
rlabel metal2 373352 2702 373352 2702 0 la_data_in[28]
rlabel metal2 378840 4102 378840 4102 0 la_data_in[29]
rlabel metal3 202944 55496 202944 55496 0 la_data_in[2]
rlabel metal2 383768 392 383768 392 0 la_data_in[30]
rlabel metal3 312704 55832 312704 55832 0 la_data_in[31]
rlabel metal3 312984 59416 312984 59416 0 la_data_in[32]
rlabel metal2 401688 4158 401688 4158 0 la_data_in[33]
rlabel metal2 406952 392 406952 392 0 la_data_in[34]
rlabel metal3 367948 7672 367948 7672 0 la_data_in[35]
rlabel metal2 418600 392 418600 392 0 la_data_in[36]
rlabel metal2 423976 392 423976 392 0 la_data_in[37]
rlabel metal3 428904 6776 428904 6776 0 la_data_in[38]
rlabel metal2 339682 60088 339682 60088 0 la_data_in[39]
rlabel metal2 230328 3150 230328 3150 0 la_data_in[3]
rlabel metal2 440944 392 440944 392 0 la_data_in[40]
rlabel metal2 447104 392 447104 392 0 la_data_in[41]
rlabel metal2 452480 392 452480 392 0 la_data_in[42]
rlabel metal2 354690 60088 354690 60088 0 la_data_in[43]
rlabel metal2 358162 60088 358162 60088 0 la_data_in[44]
rlabel metal2 361690 60088 361690 60088 0 la_data_in[45]
rlabel metal2 475664 392 475664 392 0 la_data_in[46]
rlabel metal2 481040 392 481040 392 0 la_data_in[47]
rlabel metal2 487312 11760 487312 11760 0 la_data_in[48]
rlabel metal2 376642 60088 376642 60088 0 la_data_in[49]
rlabel metal2 236040 4046 236040 4046 0 la_data_in[4]
rlabel metal2 498008 392 498008 392 0 la_data_in[50]
rlabel metal2 504224 392 504224 392 0 la_data_in[51]
rlabel metal3 386904 59416 386904 59416 0 la_data_in[52]
rlabel metal3 392784 55496 392784 55496 0 la_data_in[53]
rlabel metal2 521192 392 521192 392 0 la_data_in[54]
rlabel metal2 527352 4886 527352 4886 0 la_data_in[55]
rlabel metal1 401856 59192 401856 59192 0 la_data_in[56]
rlabel metal2 405048 39060 405048 39060 0 la_data_in[57]
rlabel metal2 544432 11760 544432 11760 0 la_data_in[58]
rlabel metal2 549752 392 549752 392 0 la_data_in[59]
rlabel metal2 241752 3318 241752 3318 0 la_data_in[5]
rlabel metal2 555128 392 555128 392 0 la_data_in[60]
rlabel metal3 560952 4984 560952 4984 0 la_data_in[61]
rlabel metal2 566720 392 566720 392 0 la_data_in[62]
rlabel metal3 571704 10136 571704 10136 0 la_data_in[63]
rlabel metal2 217434 60088 217434 60088 0 la_data_in[6]
rlabel metal3 220584 59416 220584 59416 0 la_data_in[7]
rlabel metal2 258888 3262 258888 3262 0 la_data_in[8]
rlabel metal2 264600 3990 264600 3990 0 la_data_in[9]
rlabel metal2 215096 4102 215096 4102 0 la_data_out[0]
rlabel metal2 272216 3150 272216 3150 0 la_data_out[10]
rlabel metal3 239848 56728 239848 56728 0 la_data_out[11]
rlabel metal3 243208 55496 243208 55496 0 la_data_out[12]
rlabel metal2 289128 392 289128 392 0 la_data_out[13]
rlabel metal2 295064 1470 295064 1470 0 la_data_out[14]
rlabel metal2 252266 60088 252266 60088 0 la_data_out[15]
rlabel metal2 306152 392 306152 392 0 la_data_out[16]
rlabel metal3 261688 56840 261688 56840 0 la_data_out[17]
rlabel metal1 262528 59192 262528 59192 0 la_data_out[18]
rlabel metal2 267218 60088 267218 60088 0 la_data_out[19]
rlabel metal2 220416 392 220416 392 0 la_data_out[1]
rlabel metal2 329336 5726 329336 5726 0 la_data_out[20]
rlabel metal2 334656 392 334656 392 0 la_data_out[21]
rlabel metal2 340088 392 340088 392 0 la_data_out[22]
rlabel metal2 346248 392 346248 392 0 la_data_out[23]
rlabel metal2 285698 60088 285698 60088 0 la_data_out[24]
rlabel metal2 289282 60088 289282 60088 0 la_data_out[25]
rlabel metal2 363608 3150 363608 3150 0 la_data_out[26]
rlabel metal2 368592 392 368592 392 0 la_data_out[27]
rlabel metal2 374808 392 374808 392 0 la_data_out[28]
rlabel metal2 380240 392 380240 392 0 la_data_out[29]
rlabel metal3 207088 56504 207088 56504 0 la_data_out[2]
rlabel metal2 307706 60088 307706 60088 0 la_data_out[30]
rlabel metal2 311234 60088 311234 60088 0 la_data_out[31]
rlabel metal2 314762 60088 314762 60088 0 la_data_out[32]
rlabel metal2 403368 392 403368 392 0 la_data_out[33]
rlabel metal2 408800 392 408800 392 0 la_data_out[34]
rlabel metal2 330120 33040 330120 33040 0 la_data_out[35]
rlabel metal2 329392 11760 329392 11760 0 la_data_out[36]
rlabel metal2 425712 392 425712 392 0 la_data_out[37]
rlabel metal2 432152 5726 432152 5726 0 la_data_out[38]
rlabel metal2 437304 392 437304 392 0 la_data_out[39]
rlabel metal3 207984 55496 207984 55496 0 la_data_out[3]
rlabel metal2 355320 37296 355320 37296 0 la_data_out[40]
rlabel metal2 448896 392 448896 392 0 la_data_out[41]
rlabel metal2 454272 392 454272 392 0 la_data_out[42]
rlabel metal1 354928 59192 354928 59192 0 la_data_out[43]
rlabel metal2 359688 55762 359688 55762 0 la_data_out[44]
rlabel metal2 363146 60088 363146 60088 0 la_data_out[45]
rlabel metal2 477456 392 477456 392 0 la_data_out[46]
rlabel metal2 482832 392 482832 392 0 la_data_out[47]
rlabel metal2 489272 3990 489272 3990 0 la_data_out[48]
rlabel metal2 494424 392 494424 392 0 la_data_out[49]
rlabel metal2 237944 3262 237944 3262 0 la_data_out[4]
rlabel metal3 382648 55496 382648 55496 0 la_data_out[50]
rlabel metal2 385154 60088 385154 60088 0 la_data_out[51]
rlabel metal2 512344 2702 512344 2702 0 la_data_out[52]
rlabel metal2 517832 5670 517832 5670 0 la_data_out[53]
rlabel metal2 522984 392 522984 392 0 la_data_out[54]
rlabel metal2 400106 60088 400106 60088 0 la_data_out[55]
rlabel metal2 403634 60088 403634 60088 0 la_data_out[56]
rlabel metal2 407218 60088 407218 60088 0 la_data_out[57]
rlabel metal2 546392 3150 546392 3150 0 la_data_out[58]
rlabel metal2 551544 392 551544 392 0 la_data_out[59]
rlabel metal2 215306 60088 215306 60088 0 la_data_out[5]
rlabel metal3 488096 26040 488096 26040 0 la_data_out[60]
rlabel metal2 563136 392 563136 392 0 la_data_out[61]
rlabel metal2 568512 392 568512 392 0 la_data_out[62]
rlabel metal2 574728 392 574728 392 0 la_data_out[63]
rlabel metal2 218834 60088 218834 60088 0 la_data_out[6]
rlabel metal2 222362 60088 222362 60088 0 la_data_out[7]
rlabel metal2 260792 5670 260792 5670 0 la_data_out[8]
rlabel metal2 265944 392 265944 392 0 la_data_out[9]
rlabel metal3 216440 4984 216440 4984 0 la_oenb[0]
rlabel metal2 235256 34650 235256 34650 0 la_oenb[10]
rlabel metal2 238826 60088 238826 60088 0 la_oenb[11]
rlabel metal2 242298 60088 242298 60088 0 la_oenb[12]
rlabel metal2 291256 2366 291256 2366 0 la_oenb[13]
rlabel metal2 266280 32144 266280 32144 0 la_oenb[14]
rlabel metal2 302680 2310 302680 2310 0 la_oenb[15]
rlabel metal2 308392 2646 308392 2646 0 la_oenb[16]
rlabel metal2 314216 3318 314216 3318 0 la_oenb[17]
rlabel metal2 264306 60088 264306 60088 0 la_oenb[18]
rlabel metal2 267288 57652 267288 57652 0 la_oenb[19]
rlabel metal2 222712 2478 222712 2478 0 la_oenb[1]
rlabel metal2 331240 2534 331240 2534 0 la_oenb[20]
rlabel metal2 336952 2478 336952 2478 0 la_oenb[21]
rlabel metal3 310856 54712 310856 54712 0 la_oenb[22]
rlabel metal2 282786 60088 282786 60088 0 la_oenb[23]
rlabel metal2 353416 392 353416 392 0 la_oenb[24]
rlabel metal2 359688 11760 359688 11760 0 la_oenb[25]
rlabel metal3 296240 55496 296240 55496 0 la_oenb[26]
rlabel metal2 297738 60088 297738 60088 0 la_oenb[27]
rlabel metal2 376936 2366 376936 2366 0 la_oenb[28]
rlabel metal2 382648 2310 382648 2310 0 la_oenb[29]
rlabel metal2 228536 2422 228536 2422 0 la_oenb[2]
rlabel metal3 310408 55496 310408 55496 0 la_oenb[30]
rlabel metal3 313824 55496 313824 55496 0 la_oenb[31]
rlabel metal2 316218 60088 316218 60088 0 la_oenb[32]
rlabel metal2 405496 5782 405496 5782 0 la_oenb[33]
rlabel metal2 410592 392 410592 392 0 la_oenb[34]
rlabel metal3 416360 4984 416360 4984 0 la_oenb[35]
rlabel metal3 332248 55496 332248 55496 0 la_oenb[36]
rlabel metal2 334698 60088 334698 60088 0 la_oenb[37]
rlabel metal2 433776 392 433776 392 0 la_oenb[38]
rlabel metal2 439768 3262 439768 3262 0 la_oenb[39]
rlabel metal2 234136 2366 234136 2366 0 la_oenb[3]
rlabel metal2 445368 11760 445368 11760 0 la_oenb[40]
rlabel metal2 450688 392 450688 392 0 la_oenb[41]
rlabel metal3 456568 4984 456568 4984 0 la_oenb[42]
rlabel metal2 356706 60088 356706 60088 0 la_oenb[43]
rlabel metal1 359912 59416 359912 59416 0 la_oenb[44]
rlabel metal2 474040 3206 474040 3206 0 la_oenb[45]
rlabel metal2 479248 392 479248 392 0 la_oenb[46]
rlabel metal3 428456 31192 428456 31192 0 la_oenb[47]
rlabel metal2 490840 392 490840 392 0 la_oenb[48]
rlabel metal2 496888 4830 496888 4830 0 la_oenb[49]
rlabel metal2 239848 2310 239848 2310 0 la_oenb[4]
rlabel metal2 502488 11760 502488 11760 0 la_oenb[50]
rlabel metal2 386666 60088 386666 60088 0 la_oenb[51]
rlabel metal3 452032 47880 452032 47880 0 la_oenb[52]
rlabel metal2 519736 4046 519736 4046 0 la_oenb[53]
rlabel metal3 524384 4984 524384 4984 0 la_oenb[54]
rlabel metal3 404544 55496 404544 55496 0 la_oenb[55]
rlabel metal2 405090 60088 405090 60088 0 la_oenb[56]
rlabel metal2 542696 2534 542696 2534 0 la_oenb[57]
rlabel metal2 548296 2478 548296 2478 0 la_oenb[58]
rlabel metal2 553336 392 553336 392 0 la_oenb[59]
rlabel metal2 245560 4886 245560 4886 0 la_oenb[5]
rlabel metal2 559720 2422 559720 2422 0 la_oenb[60]
rlabel metal2 565432 2366 565432 2366 0 la_oenb[61]
rlabel metal2 427098 60088 427098 60088 0 la_oenb[62]
rlabel metal2 430626 60088 430626 60088 0 la_oenb[63]
rlabel metal2 220346 60088 220346 60088 0 la_oenb[6]
rlabel metal2 257096 2534 257096 2534 0 la_oenb[7]
rlabel metal2 262696 2478 262696 2478 0 la_oenb[8]
rlabel metal2 268408 2422 268408 2422 0 la_oenb[9]
rlabel metal2 432082 60088 432082 60088 0 user_irq[0]
rlabel metal2 433608 37170 433608 37170 0 user_irq[1]
rlabel metal3 433832 59416 433832 59416 0 user_irq[2]
rlabel metal2 10696 392 10696 392 0 wb_clk_i
rlabel metal2 13384 3150 13384 3150 0 wb_rst_i
rlabel metal2 15176 18270 15176 18270 0 wbs_ack_o
rlabel metal2 72450 60088 72450 60088 0 wbs_adr_i[0]
rlabel metal2 87752 3150 87752 3150 0 wbs_adr_i[10]
rlabel metal2 117922 60088 117922 60088 0 wbs_adr_i[11]
rlabel metal2 99064 4046 99064 4046 0 wbs_adr_i[12]
rlabel metal2 104552 11760 104552 11760 0 wbs_adr_i[13]
rlabel metal2 127848 32452 127848 32452 0 wbs_adr_i[14]
rlabel metal2 128520 36176 128520 36176 0 wbs_adr_i[15]
rlabel metal2 122024 3990 122024 3990 0 wbs_adr_i[16]
rlabel metal2 127624 3206 127624 3206 0 wbs_adr_i[17]
rlabel metal3 143136 59416 143136 59416 0 wbs_adr_i[18]
rlabel metal3 146664 59416 146664 59416 0 wbs_adr_i[19]
rlabel metal2 30352 11760 30352 11760 0 wbs_adr_i[1]
rlabel metal2 144592 5880 144592 5880 0 wbs_adr_i[20]
rlabel metal2 150584 2366 150584 2366 0 wbs_adr_i[21]
rlabel metal2 156184 2646 156184 2646 0 wbs_adr_i[22]
rlabel metal2 161504 392 161504 392 0 wbs_adr_i[23]
rlabel metal2 166936 392 166936 392 0 wbs_adr_i[24]
rlabel metal3 171472 4984 171472 4984 0 wbs_adr_i[25]
rlabel metal2 173362 60088 173362 60088 0 wbs_adr_i[26]
rlabel metal3 181776 4872 181776 4872 0 wbs_adr_i[27]
rlabel metal2 190344 3150 190344 3150 0 wbs_adr_i[28]
rlabel metal2 196056 3318 196056 3318 0 wbs_adr_i[29]
rlabel metal2 37464 392 37464 392 0 wbs_adr_i[2]
rlabel metal2 188314 60088 188314 60088 0 wbs_adr_i[30]
rlabel metal2 191842 60088 191842 60088 0 wbs_adr_i[31]
rlabel metal2 45528 11760 45528 11760 0 wbs_adr_i[3]
rlabel metal2 52640 392 52640 392 0 wbs_adr_i[4]
rlabel metal2 95914 60088 95914 60088 0 wbs_adr_i[5]
rlabel metal2 99442 60088 99442 60088 0 wbs_adr_i[6]
rlabel metal2 102970 60088 102970 60088 0 wbs_adr_i[7]
rlabel metal2 75824 392 75824 392 0 wbs_adr_i[8]
rlabel metal2 82040 4102 82040 4102 0 wbs_adr_i[9]
rlabel metal2 17304 2702 17304 2702 0 wbs_cyc_i
rlabel metal2 24920 2702 24920 2702 0 wbs_dat_i[0]
rlabel metal2 89656 5670 89656 5670 0 wbs_dat_i[10]
rlabel metal2 95368 3990 95368 3990 0 wbs_dat_i[11]
rlabel metal2 101080 2534 101080 2534 0 wbs_dat_i[12]
rlabel metal2 126434 60088 126434 60088 0 wbs_dat_i[13]
rlabel metal2 112504 2366 112504 2366 0 wbs_dat_i[14]
rlabel metal2 118216 2590 118216 2590 0 wbs_dat_i[15]
rlabel metal2 123928 3150 123928 3150 0 wbs_dat_i[16]
rlabel metal2 141386 60088 141386 60088 0 wbs_dat_i[17]
rlabel metal2 142744 6104 142744 6104 0 wbs_dat_i[18]
rlabel metal2 148442 60088 148442 60088 0 wbs_dat_i[19]
rlabel metal2 32088 392 32088 392 0 wbs_dat_i[1]
rlabel metal2 146776 2702 146776 2702 0 wbs_dat_i[20]
rlabel metal2 152488 3990 152488 3990 0 wbs_dat_i[21]
rlabel metal2 158200 2702 158200 2702 0 wbs_dat_i[22]
rlabel metal2 163296 392 163296 392 0 wbs_dat_i[23]
rlabel metal3 167888 4984 167888 4984 0 wbs_dat_i[24]
rlabel metal3 172536 4872 172536 4872 0 wbs_dat_i[25]
rlabel metal2 174818 60088 174818 60088 0 wbs_dat_i[26]
rlabel metal3 182336 4200 182336 4200 0 wbs_dat_i[27]
rlabel metal2 192248 3990 192248 3990 0 wbs_dat_i[28]
rlabel metal3 194320 6328 194320 6328 0 wbs_dat_i[29]
rlabel metal2 40152 2702 40152 2702 0 wbs_dat_i[2]
rlabel metal2 188496 11760 188496 11760 0 wbs_dat_i[30]
rlabel metal2 193438 60088 193438 60088 0 wbs_dat_i[31]
rlabel metal2 47264 392 47264 392 0 wbs_dat_i[3]
rlabel metal2 54432 392 54432 392 0 wbs_dat_i[4]
rlabel metal2 95928 57652 95928 57652 0 wbs_dat_i[5]
rlabel metal2 100898 60088 100898 60088 0 wbs_dat_i[6]
rlabel metal2 72520 6510 72520 6510 0 wbs_dat_i[7]
rlabel metal2 77616 392 77616 392 0 wbs_dat_i[8]
rlabel metal2 82992 392 82992 392 0 wbs_dat_i[9]
rlabel metal2 26824 2646 26824 2646 0 wbs_dat_o[0]
rlabel metal2 94920 31192 94920 31192 0 wbs_dat_o[10]
rlabel metal2 97272 2478 97272 2478 0 wbs_dat_o[11]
rlabel metal2 102760 7350 102760 7350 0 wbs_dat_o[12]
rlabel metal2 127890 60088 127890 60088 0 wbs_dat_o[13]
rlabel metal2 114408 2422 114408 2422 0 wbs_dat_o[14]
rlabel metal2 120120 4830 120120 4830 0 wbs_dat_o[15]
rlabel metal2 125832 3150 125832 3150 0 wbs_dat_o[16]
rlabel metal2 143094 60088 143094 60088 0 wbs_dat_o[17]
rlabel metal2 146426 60088 146426 60088 0 wbs_dat_o[18]
rlabel metal2 142968 3598 142968 3598 0 wbs_dat_o[19]
rlabel metal2 34440 2478 34440 2478 0 wbs_dat_o[1]
rlabel metal2 148680 2310 148680 2310 0 wbs_dat_o[20]
rlabel metal2 154392 2702 154392 2702 0 wbs_dat_o[21]
rlabel metal2 160104 2702 160104 2702 0 wbs_dat_o[22]
rlabel metal2 165088 392 165088 392 0 wbs_dat_o[23]
rlabel metal3 169736 55496 169736 55496 0 wbs_dat_o[24]
rlabel metal2 172018 60088 172018 60088 0 wbs_dat_o[25]
rlabel metal2 174888 57540 174888 57540 0 wbs_dat_o[26]
rlabel metal2 188440 2366 188440 2366 0 wbs_dat_o[27]
rlabel metal2 194152 2702 194152 2702 0 wbs_dat_o[28]
rlabel metal2 199976 2478 199976 2478 0 wbs_dat_o[29]
rlabel metal2 41048 392 41048 392 0 wbs_dat_o[2]
rlabel metal2 190386 60088 190386 60088 0 wbs_dat_o[30]
rlabel metal3 193592 59416 193592 59416 0 wbs_dat_o[31]
rlabel metal2 49056 392 49056 392 0 wbs_dat_o[3]
rlabel metal2 57288 2534 57288 2534 0 wbs_dat_o[4]
rlabel metal2 97986 60088 97986 60088 0 wbs_dat_o[5]
rlabel metal2 100968 31836 100968 31836 0 wbs_dat_o[6]
rlabel metal2 74424 2310 74424 2310 0 wbs_dat_o[7]
rlabel metal2 80136 2366 80136 2366 0 wbs_dat_o[8]
rlabel metal2 85848 2422 85848 2422 0 wbs_dat_o[9]
rlabel metal2 28616 28350 28616 28350 0 wbs_sel_i[0]
rlabel metal2 80962 60088 80962 60088 0 wbs_sel_i[1]
rlabel metal2 43960 2422 43960 2422 0 wbs_sel_i[2]
rlabel metal2 51576 2478 51576 2478 0 wbs_sel_i[3]
rlabel metal2 19208 2310 19208 2310 0 wbs_stb_i
rlabel metal2 70994 60088 70994 60088 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
